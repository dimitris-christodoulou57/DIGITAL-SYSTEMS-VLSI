magic
tech scmos
timestamp 1544468751
<< pwell >>
rect -14 -22 37 -4
rect 71 -23 137 -5
rect 154 -17 166 -4
rect 66 -67 78 -54
<< nwell >>
rect -13 7 35 28
rect 72 6 136 27
rect 153 4 167 17
rect 65 -46 79 -33
<< polysilicon >>
rect -6 14 -4 21
rect 2 14 4 21
rect 10 14 12 21
rect 18 14 20 21
rect 26 14 28 21
rect 79 14 81 21
rect 87 14 89 21
rect 95 14 97 21
rect 103 14 105 21
rect 111 14 113 21
rect 119 14 121 21
rect 127 14 129 21
rect -6 -10 -4 11
rect 2 -10 4 11
rect 10 -10 12 11
rect 18 -10 20 11
rect 26 -10 28 11
rect 79 -10 81 11
rect 87 -10 89 11
rect 95 -10 97 11
rect 103 -10 105 11
rect 111 -10 113 11
rect 119 -10 121 11
rect 127 -10 129 11
rect 159 8 161 10
rect 159 -5 161 5
rect -6 -22 -4 -13
rect 2 -22 4 -13
rect 10 -22 12 -13
rect 18 -22 20 -13
rect 26 -22 28 -13
rect 79 -22 81 -13
rect 87 -22 89 -13
rect 95 -22 97 -13
rect 103 -28 105 -13
rect 111 -22 113 -13
rect 119 -22 121 -13
rect 127 -22 129 -13
rect 159 -16 161 -8
rect 71 -42 73 -40
rect 71 -55 73 -45
rect 71 -66 73 -58
<< ndiffusion >>
rect 158 -8 159 -5
rect 161 -8 162 -5
rect -7 -13 -6 -10
rect -4 -13 2 -10
rect 4 -13 5 -10
rect 9 -13 10 -10
rect 12 -13 13 -10
rect 17 -13 18 -10
rect 20 -13 21 -10
rect 25 -13 26 -10
rect 28 -13 29 -10
rect 78 -13 79 -10
rect 81 -13 82 -10
rect 86 -13 87 -10
rect 89 -13 90 -10
rect 94 -13 95 -10
rect 97 -13 98 -10
rect 102 -13 103 -10
rect 105 -13 106 -10
rect 110 -13 111 -10
rect 113 -13 119 -10
rect 121 -13 127 -10
rect 129 -13 130 -10
rect 70 -58 71 -55
rect 73 -58 74 -55
<< pdiffusion >>
rect -7 11 -6 14
rect -4 11 -3 14
rect 1 11 2 14
rect 4 11 5 14
rect 9 11 10 14
rect 12 11 13 14
rect 17 11 18 14
rect 20 11 26 14
rect 28 11 29 14
rect 78 11 79 14
rect 81 11 87 14
rect 89 11 95 14
rect 97 11 98 14
rect 102 11 103 14
rect 105 11 106 14
rect 110 11 111 14
rect 113 11 114 14
rect 118 11 119 14
rect 121 11 122 14
rect 126 11 127 14
rect 129 11 130 14
rect 158 5 159 8
rect 161 5 162 8
rect 70 -45 71 -42
rect 73 -45 74 -42
<< metal1 >>
rect -13 24 13 27
rect 17 24 35 27
rect 72 24 98 27
rect -11 18 8 21
rect -11 15 -8 18
rect 5 15 8 18
rect 14 15 17 24
rect 102 24 136 27
rect 99 15 102 23
rect -3 2 0 11
rect 5 8 8 11
rect 30 8 33 11
rect 5 5 33 8
rect 106 18 126 21
rect 106 15 109 18
rect 123 15 126 18
rect 74 8 77 11
rect 107 8 110 11
rect 74 5 110 8
rect 115 2 118 11
rect 131 2 134 11
rect 158 13 166 16
rect 154 9 157 13
rect 163 2 166 5
rect -13 -1 54 2
rect 72 -1 155 2
rect 5 -10 8 -1
rect 13 -7 33 -4
rect 13 -10 16 -7
rect 30 -10 33 -7
rect -11 -18 -8 -14
rect 22 -18 25 -14
rect -13 -22 -12 -19
rect -8 -22 21 -19
rect 25 -22 35 -19
rect 51 -25 54 -1
rect 82 -7 102 -4
rect 82 -10 85 -7
rect 99 -10 102 -7
rect 106 -10 109 -1
rect 163 -1 175 2
rect 163 -5 166 -1
rect 74 -18 77 -14
rect 91 -18 94 -14
rect 72 -22 73 -19
rect 77 -22 90 -19
rect 131 -18 134 -14
rect 154 -13 157 -9
rect 158 -16 166 -13
rect 94 -22 131 -19
rect 135 -22 136 -19
rect 51 -28 99 -25
rect 51 -49 54 -28
rect 70 -37 78 -34
rect 66 -41 69 -37
rect 75 -48 78 -45
rect 51 -52 67 -49
rect 75 -51 86 -48
rect 75 -55 78 -51
rect 66 -63 69 -59
rect 70 -66 78 -63
<< ntransistor >>
rect 159 -8 161 -5
rect -6 -13 -4 -10
rect 2 -13 4 -10
rect 10 -13 12 -10
rect 18 -13 20 -10
rect 26 -13 28 -10
rect 79 -13 81 -10
rect 87 -13 89 -10
rect 95 -13 97 -10
rect 103 -13 105 -10
rect 111 -13 113 -10
rect 119 -13 121 -10
rect 127 -13 129 -10
rect 71 -58 73 -55
<< ptransistor >>
rect -6 11 -4 14
rect 2 11 4 14
rect 10 11 12 14
rect 18 11 20 14
rect 26 11 28 14
rect 79 11 81 14
rect 87 11 89 14
rect 95 11 97 14
rect 103 11 105 14
rect 111 11 113 14
rect 119 11 121 14
rect 127 11 129 14
rect 159 5 161 8
rect 71 -45 73 -42
<< polycontact >>
rect 155 -2 159 2
rect 99 -29 103 -25
rect 67 -52 71 -48
<< ndcontact >>
rect 154 -9 158 -5
rect -11 -14 -7 -10
rect 5 -14 9 -10
rect 13 -14 17 -10
rect 21 -14 25 -10
rect 29 -14 33 -10
rect 74 -14 78 -10
rect 82 -14 86 -10
rect 90 -14 94 -10
rect 98 -14 102 -10
rect 106 -14 110 -10
rect 130 -14 134 -10
rect 162 -9 166 -5
rect 66 -59 70 -55
rect 74 -59 78 -55
<< pdcontact >>
rect -11 11 -7 15
rect -3 11 1 15
rect 5 11 9 15
rect 13 11 17 15
rect 29 11 33 15
rect 74 11 78 15
rect 98 11 102 15
rect 106 11 110 15
rect 114 11 118 15
rect 122 11 126 15
rect 130 11 134 15
rect 154 5 158 9
rect 162 5 166 9
rect 66 -45 70 -41
rect 74 -45 78 -41
<< psubstratepcontact >>
rect -12 -22 -8 -18
rect 21 -22 25 -18
rect 73 -22 77 -18
rect 90 -22 94 -18
rect 154 -17 158 -13
rect 131 -22 135 -18
rect 66 -67 70 -63
<< nsubstratencontact >>
rect 13 24 17 28
rect 98 23 102 27
rect 154 13 158 17
rect 66 -37 70 -33
<< labels >>
rlabel metal1 -13 24 35 27 1 VDD
rlabel metal1 -13 -22 35 -19 5 GND
rlabel polysilicon -6 -10 -4 11 0 Cin
rlabel polysilicon 2 -10 4 11 0 B
rlabel polysilicon 10 -10 12 11 0 A
rlabel polysilicon 18 -10 20 11 0 B
rlabel polysilicon 26 -10 28 11 0 Cin
rlabel metal1 -13 -1 35 2 3 Cout'
rlabel metal1 72 24 136 27 1 VDD
rlabel metal1 72 -22 136 -19 5 GND
rlabel polysilicon 79 -10 81 11 0 A
rlabel polysilicon 87 -10 89 11 0 B
rlabel polysilicon 95 -10 97 11 0 Cin
rlabel polysilicon 111 -10 113 11 0 A
rlabel polysilicon 119 -10 121 11 0 B
rlabel polysilicon 127 -10 129 11 0 Cin
rlabel metal1 75 -51 86 -48 3 Cout
rlabel metal1 66 -37 78 -34 1 VDD
rlabel metal1 66 -66 78 -63 5 GND
rlabel metal1 154 13 166 16 1 VDD
rlabel metal1 154 -16 166 -13 5 GND
rlabel metal1 72 -1 155 2 1 Sout'
rlabel metal1 163 -1 175 2 3 Sout
<< end >>
