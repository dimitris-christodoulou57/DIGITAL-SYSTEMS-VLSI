magic
tech scmos
timestamp 1542766022
<< polysilicon >>
rect -15 14 23 16
rect -15 6 -13 14
rect -6 10 14 12
rect -6 6 -4 10
rect 3 6 5 8
rect 12 6 14 10
rect 21 6 23 14
rect -15 -22 -13 3
rect -6 -22 -4 3
rect 3 -22 5 3
rect 12 -22 14 3
rect 21 -22 23 3
rect -15 -34 -13 -25
rect -6 -34 -4 -25
rect 3 -34 5 -25
rect 12 -34 14 -25
rect 21 -34 23 -25
<< ndiffusion >>
rect -17 -25 -15 -22
rect -13 -25 -6 -22
rect -4 -25 -2 -22
rect 2 -25 3 -22
rect 5 -25 7 -22
rect 11 -25 12 -22
rect 14 -25 16 -22
rect 20 -25 21 -22
rect 23 -25 25 -22
<< pdiffusion >>
rect -17 3 -15 6
rect -13 3 -11 6
rect -7 3 -6 6
rect -4 3 -2 6
rect 2 3 3 6
rect 5 3 7 6
rect 11 3 12 6
rect 14 3 21 6
rect 23 3 25 6
<< metal1 >>
rect -23 17 31 20
rect -11 7 -8 17
rect 25 7 28 17
rect -20 -1 -17 3
rect -2 -1 1 3
rect -20 -4 1 -1
rect 7 -8 10 3
rect -23 -11 31 -8
rect -20 -18 10 -15
rect -20 -22 -17 -18
rect 7 -22 10 -18
rect 16 -22 19 -11
rect -2 -36 1 -26
rect 7 -29 10 -26
rect 25 -29 28 -26
rect 7 -32 28 -29
rect -23 -39 31 -36
<< ntransistor >>
rect -15 -25 -13 -22
rect -6 -25 -4 -22
rect 3 -25 5 -22
rect 12 -25 14 -22
rect 21 -25 23 -22
<< ptransistor >>
rect -15 3 -13 6
rect -6 3 -4 6
rect 3 3 5 6
rect 12 3 14 6
rect 21 3 23 6
<< ndcontact >>
rect -21 -26 -17 -22
rect -2 -26 2 -22
rect 7 -26 11 -22
rect 16 -26 20 -22
rect 25 -26 29 -22
<< pdcontact >>
rect -21 3 -17 7
rect -11 3 -7 7
rect -2 3 2 7
rect 7 3 11 7
rect 25 3 29 7
<< labels >>
rlabel metal1 -23 -11 31 -8 7 vout
rlabel metal1 -23 17 31 20 7 vdd
rlabel metal1 -23 -39 31 -36 7 gnd
rlabel polysilicon 3 6 5 8 1 b
rlabel polysilicon -6 10 14 12 1 a
rlabel polysilicon -15 14 23 16 1 c
<< end >>
