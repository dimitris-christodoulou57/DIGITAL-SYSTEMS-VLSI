magic
tech scmos
timestamp 1546883516
<< pwell >>
rect -47 14 -33 27
rect 64 19 78 32
rect 6 -38 50 -20
rect 6 -112 50 -94
rect 90 -117 104 -104
rect 6 -189 50 -168
rect 6 -263 50 -242
rect 6 -337 50 -316
rect 6 -411 50 -390
rect 6 -485 50 -464
rect 6 -559 50 -538
<< nwell >>
rect -47 37 -33 50
rect 64 42 78 55
rect 6 -6 50 22
rect 6 -80 50 -52
rect 90 -94 104 -81
rect 6 -154 50 -126
rect 6 -228 50 -200
rect 6 -302 50 -274
rect 6 -376 50 -348
rect 6 -450 50 -422
rect 6 -524 50 -496
<< polysilicon >>
rect 70 46 72 48
rect -41 41 -39 43
rect -41 25 -39 38
rect -41 20 -39 22
rect 18 10 20 32
rect 28 10 30 14
rect 38 10 40 38
rect 70 30 72 43
rect 70 25 72 27
rect 18 -26 20 -2
rect 28 -26 30 -2
rect 38 -26 40 -2
rect 18 -34 20 -29
rect 18 -64 20 -45
rect 28 -64 30 -29
rect 38 -64 40 -29
rect 18 -100 20 -76
rect 28 -100 30 -76
rect 38 -100 40 -76
rect 96 -90 98 -88
rect 18 -108 20 -103
rect 28 -108 30 -103
rect 18 -138 20 -120
rect 28 -138 30 -135
rect 38 -138 40 -103
rect 96 -106 98 -93
rect 96 -111 98 -109
rect 18 -177 20 -150
rect 28 -177 30 -150
rect 38 -177 40 -150
rect 18 -183 20 -180
rect 18 -212 20 -194
rect 28 -212 30 -180
rect 38 -212 40 -180
rect 18 -251 20 -224
rect 28 -251 30 -224
rect 38 -251 40 -224
rect 18 -257 20 -254
rect 28 -257 30 -254
rect 38 -257 40 -254
rect 18 -286 20 -268
rect 28 -286 30 -283
rect 38 -286 40 -271
rect 18 -325 20 -298
rect 28 -325 30 -298
rect 38 -325 40 -298
rect 18 -331 20 -328
rect 18 -360 20 -342
rect 28 -360 30 -328
rect 38 -360 40 -328
rect 18 -399 20 -372
rect 28 -399 30 -372
rect 38 -399 40 -372
rect 18 -405 20 -402
rect 28 -405 30 -402
rect 18 -434 20 -416
rect 28 -434 30 -431
rect 38 -434 40 -402
rect 18 -473 20 -446
rect 28 -473 30 -446
rect 38 -473 40 -446
rect 18 -479 20 -476
rect 18 -508 20 -490
rect 28 -508 30 -476
rect 38 -508 40 -476
rect 18 -547 20 -520
rect 28 -547 30 -520
rect 38 -547 40 -520
rect 18 -553 20 -550
rect 28 -553 30 -550
rect 38 -567 40 -550
<< ndiffusion >>
rect -43 22 -41 25
rect -39 22 -37 25
rect 68 27 70 30
rect 72 27 74 30
rect 16 -29 18 -26
rect 20 -29 22 -26
rect 26 -29 28 -26
rect 30 -29 32 -26
rect 36 -29 38 -26
rect 40 -29 42 -26
rect 16 -103 18 -100
rect 20 -103 22 -100
rect 26 -103 28 -100
rect 30 -103 32 -100
rect 36 -103 38 -100
rect 40 -103 42 -100
rect 94 -109 96 -106
rect 98 -109 100 -106
rect 16 -180 18 -177
rect 20 -180 22 -177
rect 26 -180 28 -177
rect 30 -180 32 -177
rect 36 -180 38 -177
rect 40 -180 42 -177
rect 16 -254 18 -251
rect 20 -254 22 -251
rect 26 -254 28 -251
rect 30 -254 32 -251
rect 36 -254 38 -251
rect 40 -254 42 -251
rect 16 -328 18 -325
rect 20 -328 22 -325
rect 26 -328 28 -325
rect 30 -328 32 -325
rect 36 -328 38 -325
rect 40 -328 42 -325
rect 16 -402 18 -399
rect 20 -402 22 -399
rect 26 -402 28 -399
rect 30 -402 32 -399
rect 36 -402 38 -399
rect 40 -402 42 -399
rect 17 -476 18 -473
rect 20 -476 22 -473
rect 26 -476 28 -473
rect 30 -476 32 -473
rect 36 -476 38 -473
rect 40 -476 42 -473
rect 16 -550 18 -547
rect 20 -550 22 -547
rect 26 -550 28 -547
rect 30 -550 32 -547
rect 36 -550 38 -547
rect 40 -550 42 -547
<< pdiffusion >>
rect 68 43 70 46
rect 72 43 74 46
rect -43 38 -41 41
rect -39 38 -37 41
rect 16 -2 18 10
rect 20 -2 28 10
rect 30 -2 38 10
rect 40 -2 42 10
rect 16 -76 18 -64
rect 20 -76 28 -64
rect 30 -76 38 -64
rect 40 -76 42 -64
rect 94 -93 96 -90
rect 98 -93 100 -90
rect 16 -150 18 -138
rect 20 -150 28 -138
rect 30 -150 38 -138
rect 40 -150 42 -138
rect 16 -224 18 -212
rect 20 -224 28 -212
rect 30 -224 38 -212
rect 40 -224 42 -212
rect 16 -298 18 -286
rect 20 -298 28 -286
rect 30 -298 38 -286
rect 40 -298 42 -286
rect 16 -372 18 -360
rect 20 -372 28 -360
rect 30 -372 38 -360
rect 40 -372 42 -360
rect 16 -446 18 -434
rect 20 -446 28 -434
rect 30 -446 38 -434
rect 40 -446 42 -434
rect 16 -520 18 -508
rect 20 -520 28 -508
rect 30 -520 38 -508
rect 40 -520 42 -508
<< metal1 >>
rect 64 51 78 54
rect -47 46 -33 49
rect 75 47 78 51
rect -47 42 -44 46
rect 64 38 67 43
rect -58 30 -45 33
rect -36 32 -33 38
rect 44 35 67 38
rect 76 36 121 39
rect -36 29 14 32
rect -36 25 -33 29
rect -47 18 -44 21
rect -47 15 -33 18
rect -29 -120 -26 29
rect 64 30 67 35
rect 75 23 78 26
rect 6 18 50 21
rect 64 20 78 23
rect 42 10 46 18
rect 12 -11 16 -2
rect 12 -14 54 -11
rect 22 -25 25 -14
rect 43 -25 46 -14
rect 12 -35 15 -29
rect 33 -35 36 -29
rect 6 -38 50 -35
rect -1 -48 14 -45
rect 34 -46 74 -43
rect 6 -56 50 -53
rect 42 -64 46 -56
rect 12 -85 16 -76
rect 12 -88 49 -85
rect 22 -99 25 -88
rect 43 -99 46 -88
rect 71 -97 74 -46
rect 90 -85 104 -82
rect 101 -89 104 -85
rect 90 -97 93 -93
rect 71 -100 93 -97
rect 12 -109 15 -103
rect 33 -109 36 -103
rect 6 -112 50 -109
rect -29 -123 14 -120
rect -29 -268 -26 -123
rect 6 -130 50 -127
rect 42 -138 46 -130
rect 12 -159 16 -150
rect 12 -162 49 -159
rect 22 -176 25 -162
rect 43 -176 46 -162
rect 12 -186 15 -180
rect 33 -186 36 -180
rect 6 -189 50 -186
rect -1 -197 14 -194
rect 34 -196 65 -193
rect 6 -204 50 -201
rect 42 -212 46 -204
rect 12 -233 16 -224
rect 12 -236 49 -233
rect 22 -250 25 -236
rect 43 -250 46 -236
rect 12 -260 15 -254
rect 33 -260 36 -254
rect 6 -263 50 -260
rect -29 -271 14 -268
rect -29 -416 -26 -271
rect 6 -278 50 -275
rect 42 -286 46 -278
rect 12 -307 16 -298
rect 12 -310 49 -307
rect 22 -324 25 -310
rect 43 -324 46 -310
rect 12 -334 15 -328
rect 33 -334 36 -328
rect 6 -337 50 -334
rect 71 -341 74 -100
rect 90 -106 93 -100
rect 102 -100 111 -97
rect 101 -113 104 -110
rect 90 -116 104 -113
rect -1 -345 14 -342
rect 34 -344 74 -341
rect 6 -352 50 -349
rect 42 -360 46 -352
rect 12 -381 16 -372
rect 12 -384 49 -381
rect 22 -398 25 -384
rect 43 -398 46 -384
rect 12 -408 15 -402
rect 33 -408 36 -402
rect 6 -411 50 -408
rect -29 -419 14 -416
rect 6 -426 50 -423
rect 42 -434 46 -426
rect 12 -455 16 -446
rect 12 -458 49 -455
rect 22 -472 25 -458
rect 43 -472 46 -458
rect 13 -482 16 -476
rect 33 -482 36 -476
rect 6 -485 50 -482
rect -1 -493 14 -490
rect 34 -491 65 -488
rect 6 -500 50 -497
rect 42 -508 46 -500
rect 12 -529 16 -520
rect 12 -532 49 -529
rect 22 -546 25 -532
rect 43 -546 46 -532
rect 12 -556 15 -550
rect 33 -556 36 -550
rect 6 -559 50 -556
rect 118 -564 121 36
rect 44 -567 121 -564
<< ntransistor >>
rect -41 22 -39 25
rect 70 27 72 30
rect 18 -29 20 -26
rect 28 -29 30 -26
rect 38 -29 40 -26
rect 18 -103 20 -100
rect 28 -103 30 -100
rect 38 -103 40 -100
rect 96 -109 98 -106
rect 18 -180 20 -177
rect 28 -180 30 -177
rect 38 -180 40 -177
rect 18 -254 20 -251
rect 28 -254 30 -251
rect 38 -254 40 -251
rect 18 -328 20 -325
rect 28 -328 30 -325
rect 38 -328 40 -325
rect 18 -402 20 -399
rect 28 -402 30 -399
rect 38 -402 40 -399
rect 18 -476 20 -473
rect 28 -476 30 -473
rect 38 -476 40 -473
rect 18 -550 20 -547
rect 28 -550 30 -547
rect 38 -550 40 -547
<< ptransistor >>
rect 70 43 72 46
rect -41 38 -39 41
rect 18 -2 20 10
rect 28 -2 30 10
rect 38 -2 40 10
rect 18 -76 20 -64
rect 28 -76 30 -64
rect 38 -76 40 -64
rect 96 -93 98 -90
rect 18 -150 20 -138
rect 28 -150 30 -138
rect 38 -150 40 -138
rect 18 -224 20 -212
rect 28 -224 30 -212
rect 38 -224 40 -212
rect 18 -298 20 -286
rect 28 -298 30 -286
rect 38 -298 40 -286
rect 18 -372 20 -360
rect 28 -372 30 -360
rect 38 -372 40 -360
rect 18 -446 20 -434
rect 28 -446 30 -434
rect 38 -446 40 -434
rect 18 -520 20 -508
rect 28 -520 30 -508
rect 38 -520 40 -508
<< polycontact >>
rect -45 29 -41 33
rect 14 28 18 32
rect 40 34 44 38
rect 72 35 76 39
rect 14 -49 18 -45
rect 30 -47 34 -43
rect 14 -124 18 -120
rect 98 -101 102 -97
rect 14 -198 18 -194
rect 30 -197 34 -193
rect 14 -272 18 -268
rect 14 -346 18 -342
rect 30 -345 34 -341
rect 14 -420 18 -416
rect 14 -494 18 -490
rect 30 -492 34 -488
rect 40 -567 44 -563
<< ndcontact >>
rect -47 21 -43 25
rect -37 21 -33 25
rect 64 26 68 30
rect 74 26 78 30
rect 12 -29 16 -25
rect 22 -29 26 -25
rect 32 -29 36 -25
rect 42 -29 46 -25
rect 12 -103 16 -99
rect 22 -103 26 -99
rect 32 -103 36 -99
rect 42 -103 46 -99
rect 90 -110 94 -106
rect 100 -110 104 -106
rect 12 -180 16 -176
rect 22 -180 26 -176
rect 32 -180 36 -176
rect 42 -180 46 -176
rect 12 -254 16 -250
rect 22 -254 26 -250
rect 32 -254 36 -250
rect 42 -254 46 -250
rect 12 -328 16 -324
rect 22 -328 26 -324
rect 32 -328 36 -324
rect 42 -328 46 -324
rect 12 -402 16 -398
rect 22 -402 26 -398
rect 32 -402 36 -398
rect 42 -402 46 -398
rect 13 -476 17 -472
rect 22 -476 26 -472
rect 32 -476 36 -472
rect 42 -476 46 -472
rect 12 -550 16 -546
rect 22 -550 26 -546
rect 32 -550 36 -546
rect 42 -550 46 -546
<< pdcontact >>
rect 64 43 68 47
rect 74 43 78 47
rect -47 38 -43 42
rect -37 38 -33 42
rect 12 -2 16 10
rect 42 -2 46 10
rect 12 -76 16 -64
rect 42 -76 46 -64
rect 90 -93 94 -89
rect 100 -93 104 -89
rect 12 -150 16 -138
rect 42 -150 46 -138
rect 12 -224 16 -212
rect 42 -224 46 -212
rect 12 -298 16 -286
rect 42 -298 46 -286
rect 12 -372 16 -360
rect 42 -372 46 -360
rect 12 -446 16 -434
rect 42 -446 46 -434
rect 12 -520 16 -508
rect 42 -520 46 -508
<< labels >>
rlabel metal1 6 -38 50 -35 5 GND
rlabel metal1 6 18 50 21 1 VDD
rlabel metal1 6 -56 50 -53 1 VDD
rlabel metal1 6 -130 50 -127 1 VDD
rlabel metal1 6 -204 50 -201 1 VDD
rlabel metal1 6 -278 50 -275 1 VDD
rlabel metal1 6 -352 50 -349 1 VDD
rlabel metal1 6 -426 50 -423 1 VDD
rlabel metal1 6 -500 50 -497 1 VDD
rlabel metal1 6 -559 50 -556 5 GND
rlabel metal1 6 -485 50 -482 5 GND
rlabel metal1 6 -411 50 -408 5 GND
rlabel metal1 6 -337 50 -334 5 GND
rlabel metal1 6 -263 50 -260 5 GND
rlabel metal1 6 -189 50 -186 5 GND
rlabel metal1 6 -112 50 -109 5 GND
rlabel metal1 -47 46 -33 49 1 VDD
rlabel metal1 -47 15 -33 18 5 GND
rlabel metal1 64 51 78 54 1 VDD
rlabel metal1 64 20 78 23 5 GND
rlabel metal1 44 35 67 38 5 A2
rlabel metal1 44 35 67 38 5 A2'
rlabel metal1 118 -278 121 39 3 A2
rlabel metal1 -58 30 -43 33 5 A0
rlabel metal1 -36 29 -23 32 1 A0'
rlabel metal1 -1 -493 16 -490 1 A0
rlabel metal1 -1 -345 16 -342 1 A0
rlabel metal1 -1 -197 16 -194 1 A0
rlabel metal1 -1 -48 16 -45 1 A0
rlabel metal1 32 -196 65 -193 1 A1
rlabel metal1 32 -491 65 -488 1 A1
rlabel metal1 71 -100 93 -97 1 A1'
rlabel metal1 100 -100 111 -97 1 A1
rlabel metal1 90 -116 104 -113 5 GND
rlabel metal1 90 -85 104 -82 1 VDD
rlabel metal1 12 -14 54 -11 3 Z0
rlabel metal1 12 -88 49 -85 3 Z1
rlabel metal1 12 -162 49 -159 3 z2
rlabel metal1 12 -236 49 -233 3 Z3
rlabel metal1 12 -310 49 -307 3 Z4
rlabel metal1 12 -384 49 -381 3 Z5
rlabel metal1 12 -458 49 -455 3 Z6
rlabel metal1 12 -532 49 -529 3 Z7
<< end >>
