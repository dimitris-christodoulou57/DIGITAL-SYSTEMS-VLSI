* SPICE3 file created from inverter.ext - technology: scmos

.include 0.25-models

M1000 out in vdd vdd CMOSP w=3u l=2u
+  ad=19p pd=18u as=19p ps=18u
M1001 out in gnd gnd CMOSN w=3u l=2u
+  ad=19p pd=18u as=19p ps=18u
C0 gnd in 2.48fF
C1 vdd in 2.97fF

vvdd vdd 0 2.5v DC

vin in 0 pwl
+0ns 0v
+2.8ns 0v
+3ns 2.5v
+8.8ns 2.5v
+9ns 0v
+14.8ns 0v
+15ns 2.5v
+20.8ns 2.5v
+21ns 0v

.tran 10ps 25ns

*Inertial Delay UP
.meas tran t1 trig v(in) val=1.25 rise=1
+targ v(out) val=1.25 fall=1

*Inertial Delay DOWN
.meas tran t2 trig v(in) val=1.25 fall=1
+targ v(out) val=1.25 rise=1

*RISE
.meas tran rise trig v(out) val=0.25 rise=1
+targ v(out) val=2.25 rise=1

*FALL
.meas tran fall trig v(out) val=2.25 fall=1
+targ v(out) val=0.25 fall=1

.end
