magic
tech scmos
timestamp 1539623934
<< pwell >>
rect -9 -21 5 -4
<< nwell >>
rect -9 -3 5 15
<< polysilicon >>
rect -3 5 -1 7
rect -3 -8 -1 2
rect -3 -13 -1 -11
<< ndiffusion >>
rect -4 -11 -3 -8
rect -1 -11 0 -8
<< pdiffusion >>
rect -4 2 -3 5
rect -1 2 0 5
<< metal1 >>
rect -4 10 4 14
rect -8 6 -4 10
rect 0 -1 4 2
rect -15 -5 -7 -1
rect 0 -5 10 -1
rect 0 -8 4 -5
rect -8 -16 -4 -12
rect -4 -20 4 -16
<< ntransistor >>
rect -3 -11 -1 -8
<< ptransistor >>
rect -3 2 -1 5
<< polycontact >>
rect -7 -5 -3 -1
<< ndcontact >>
rect -8 -12 -4 -8
rect 0 -12 4 -8
<< pdcontact >>
rect -8 2 -4 6
rect 0 2 4 6
<< psubstratepcontact >>
rect -8 -20 -4 -16
<< nsubstratencontact >>
rect -8 10 -4 14
<< labels >>
rlabel metal1 0 -5 10 -1 3 out
rlabel metal1 -15 -5 -5 -1 7 in
rlabel metal1 -8 10 4 14 0 vdd
rlabel metal1 -8 -20 4 -16 0 gnd
<< end >>
