magic
tech scmos
timestamp 1546884218
<< pwell >>
rect 6 -38 50 -20
<< nwell >>
rect 6 -6 50 22
<< polysilicon >>
rect 18 10 20 12
rect 28 10 30 12
rect 38 10 40 12
rect 18 -26 20 -2
rect 28 -26 30 -2
rect 38 -26 40 -2
rect 18 -31 20 -29
rect 28 -31 30 -29
rect 38 -31 40 -29
<< ndiffusion >>
rect 16 -29 18 -26
rect 20 -29 22 -26
rect 26 -29 28 -26
rect 30 -29 32 -26
rect 36 -29 38 -26
rect 40 -29 42 -26
<< pdiffusion >>
rect 16 -2 18 10
rect 20 -2 28 10
rect 30 -2 38 10
rect 40 -2 42 10
<< metal1 >>
rect 6 18 50 21
rect 42 10 46 18
rect 12 -11 16 -2
rect 12 -14 54 -11
rect 22 -25 25 -14
rect 43 -25 46 -14
rect 12 -35 15 -29
rect 33 -35 36 -29
rect 6 -38 50 -35
<< ntransistor >>
rect 18 -29 20 -26
rect 28 -29 30 -26
rect 38 -29 40 -26
<< ptransistor >>
rect 18 -2 20 10
rect 28 -2 30 10
rect 38 -2 40 10
<< ndcontact >>
rect 12 -29 16 -25
rect 22 -29 26 -25
rect 32 -29 36 -25
rect 42 -29 46 -25
<< pdcontact >>
rect 12 -2 16 10
rect 42 -2 46 10
<< labels >>
rlabel metal1 6 -38 50 -35 5 GND
rlabel metal1 6 18 50 21 1 VDD
rlabel metal1 12 -14 54 -11 3 Z0
<< end >>
