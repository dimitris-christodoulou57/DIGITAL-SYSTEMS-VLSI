* SPICE3 file created from inverter.ext - technology: scmos

.include 0.25-models

M1000 out in vdd vdd CMOSP w=3u l=2u
+  ad=19p pd=18u as=19p ps=18u
M1001 out in 0 0 CMOSN w=3u l=2u
+  ad=19p pd=18u as=19p ps=18u

V1 vdd 0 0.7v DC
Vin in 0 0 DC
.dc Vin 0 0.7v 0.1

.control
	run
	plot v(out) v(in)
	plot -i(V1)
	let P = -(i(V1))*v(vdd)
	plot P
	print mean(-(i(V1)))
	print mean(P)
.endc

.end
