* SPICE3 file latch.spice

.include 0.25-models

.subckt inv drain gate source bulk
	M1 drain gate source bulk CMOSP w=18u l=3u
	M2 drain gate 0 0 CMOSN w=6u l=3u
.ends

.subckt back_inv drain gate source bulk
	M3 drain gate source bulk CMOSP w=9u l=3u
	M4 drain gate 0 0 CMOSN w=3u l=3u
.ends

Vvdd vdd 0 2.5v dc
Vclk clk 0 pwl (0 0 10ns 0 10.2ns 2.5 20ns 2.5 20.2ns 0 30ns 0 30.2ns 2.5 40ns 2.5 40.2ns 0 50ns 0 50.2ns 2.5 60ns 2.5 60.2ns 0 70ns 0 70.2ns 2.5 80 2.5 80.2ns 0)
* VDin Din 0 pwl (0 0 20ns 0 20.4ns 2.5 40ns 2.5 40.4ns 0 70ns 0 70.4ns 2.5 100ns 2.5)
VDin Din 0 pwl (0 2.5 20ns 2.5 20.4ns 0 40ns 0 40.4ns 2.5 70ns 2.5 70.4ns 0 100ns 0)

Xinv1 Dout Din vdd vdd inv
Xinv2 clk_out clk vdd vdd inv

Mclk1 Qin clk Dout vdd CMOSP w=27u l=3u
Mclk2 Qin clk_out Dout 0 CMOSN w=9u l=3u

Xinv3 Q Qin vdd vdd inv
Xinv4 Qin Q vdd vdd back_inv

.tran 10ps 110ns

.control
	run
	plot Din clk Q
