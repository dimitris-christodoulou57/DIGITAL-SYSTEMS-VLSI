magic
tech scmos
timestamp 1542765016
<< polysilicon >>
rect -16 6 -14 15
rect -5 6 -3 15
rect 6 6 8 15
rect 20 6 22 15
rect -16 -22 -14 3
rect -5 -22 -3 3
rect 6 -22 8 3
rect 20 -22 22 3
rect -16 -34 -14 -25
rect -5 -34 -3 -25
rect 6 -34 8 -25
rect 20 -34 22 -25
<< ndiffusion >>
rect -17 -25 -16 -22
rect -14 -25 -11 -22
rect -7 -25 -5 -22
rect -3 -25 0 -22
rect 4 -25 6 -22
rect 8 -25 12 -22
rect 16 -25 20 -22
rect 22 -25 25 -22
<< pdiffusion >>
rect -17 3 -16 6
rect -14 3 -5 6
rect -3 3 6 6
rect 8 3 12 6
rect 16 3 20 6
rect 22 3 25 6
<< metal1 >>
rect -23 17 31 20
rect -20 7 -17 17
rect 25 7 28 17
rect 13 -8 16 3
rect -23 -11 31 -8
rect -11 -19 16 -16
rect -11 -22 -8 -19
rect 13 -22 16 -19
rect 25 -22 28 -11
rect -20 -36 -17 -26
rect 0 -36 3 -26
rect -23 -39 31 -36
<< ntransistor >>
rect -16 -25 -14 -22
rect -5 -25 -3 -22
rect 6 -25 8 -22
rect 20 -25 22 -22
<< ptransistor >>
rect -16 3 -14 6
rect -5 3 -3 6
rect 6 3 8 6
rect 20 3 22 6
<< ndcontact >>
rect -21 -26 -17 -22
rect -11 -26 -7 -22
rect 0 -26 4 -22
rect 12 -26 16 -22
rect 25 -26 29 -22
<< pdcontact >>
rect -21 3 -17 7
rect 12 3 16 7
rect 25 3 29 7
<< labels >>
rlabel metal1 -23 -39 31 -36 7 gnd
rlabel metal1 -23 -11 31 -8 7 vout
rlabel metal1 -23 17 31 20 7 vdd
rlabel polysilicon -16 6 -14 15 1 a
rlabel polysilicon -5 6 -3 15 1 c
rlabel polysilicon 6 6 8 15 1 d
rlabel polysilicon 20 6 22 15 1 b
<< end >>
