magic
tech scmos
timestamp 1544476343
<< pwell >>
rect -1727 -8 -1676 10
rect -1642 -9 -1576 9
rect -1559 -3 -1547 10
rect -1473 -4 -1422 14
rect -1388 -5 -1322 13
rect -1305 1 -1293 14
rect -1274 -11 -1223 7
rect -1189 -12 -1123 6
rect -1106 -6 -1094 7
rect -1071 -17 -1020 1
rect -986 -18 -920 0
rect -903 -12 -891 1
rect -756 -3 -705 15
rect -671 -4 -605 14
rect -588 2 -576 15
rect -503 -12 -452 6
rect -418 -13 -352 5
rect -335 -7 -323 6
rect -260 -18 -209 0
rect -175 -19 -109 -1
rect -92 -13 -80 0
rect -14 -22 37 -4
rect 71 -23 137 -5
rect 154 -17 166 -4
rect -1647 -53 -1635 -40
rect -1393 -49 -1381 -36
rect -1194 -56 -1182 -43
rect -676 -48 -664 -35
rect -991 -62 -979 -49
rect -423 -57 -411 -44
rect -180 -63 -168 -50
rect 66 -67 78 -54
<< nwell >>
rect -1726 21 -1678 42
rect -1641 20 -1577 41
rect -1560 18 -1546 31
rect -1472 25 -1424 46
rect -1387 24 -1323 45
rect -1306 22 -1292 35
rect -1273 18 -1225 39
rect -1188 17 -1124 38
rect -1107 15 -1093 28
rect -1070 12 -1022 33
rect -985 11 -921 32
rect -755 26 -707 47
rect -670 25 -606 46
rect -589 23 -575 36
rect -904 9 -890 22
rect -502 17 -454 38
rect -417 16 -353 37
rect -1648 -32 -1634 -19
rect -1394 -28 -1380 -15
rect -336 14 -322 27
rect -259 11 -211 32
rect -174 10 -110 31
rect -93 8 -79 21
rect -13 7 35 28
rect 72 6 136 27
rect 153 4 167 17
rect -1195 -35 -1181 -22
rect -677 -27 -663 -14
rect -992 -41 -978 -28
rect -424 -36 -410 -23
rect -181 -42 -167 -29
rect 65 -46 79 -33
<< polysilicon >>
rect -1719 28 -1717 35
rect -1711 28 -1709 35
rect -1703 28 -1701 35
rect -1695 28 -1693 35
rect -1687 28 -1685 35
rect -1634 28 -1632 35
rect -1626 28 -1624 35
rect -1618 28 -1616 35
rect -1610 28 -1608 35
rect -1602 28 -1600 35
rect -1594 28 -1592 35
rect -1586 28 -1584 35
rect -1465 32 -1463 39
rect -1457 32 -1455 39
rect -1449 32 -1447 39
rect -1441 32 -1439 39
rect -1433 32 -1431 39
rect -1380 32 -1378 39
rect -1372 32 -1370 39
rect -1364 32 -1362 39
rect -1356 32 -1354 39
rect -1348 32 -1346 39
rect -1340 32 -1338 39
rect -1332 32 -1330 39
rect -1719 4 -1717 25
rect -1711 4 -1709 25
rect -1703 4 -1701 25
rect -1695 4 -1693 25
rect -1687 4 -1685 25
rect -1634 4 -1632 25
rect -1626 4 -1624 25
rect -1618 4 -1616 25
rect -1610 4 -1608 25
rect -1602 4 -1600 25
rect -1594 4 -1592 25
rect -1586 4 -1584 25
rect -1554 22 -1552 24
rect -1554 9 -1552 19
rect -1719 -8 -1717 1
rect -1711 -8 -1709 1
rect -1703 -8 -1701 1
rect -1695 -8 -1693 1
rect -1687 -8 -1685 1
rect -1634 -8 -1632 1
rect -1626 -8 -1624 1
rect -1618 -8 -1616 1
rect -1610 -14 -1608 1
rect -1602 -8 -1600 1
rect -1594 -8 -1592 1
rect -1586 -8 -1584 1
rect -1554 -2 -1552 6
rect -1465 8 -1463 29
rect -1457 8 -1455 29
rect -1449 8 -1447 29
rect -1441 8 -1439 29
rect -1433 8 -1431 29
rect -1380 8 -1378 29
rect -1372 8 -1370 29
rect -1364 8 -1362 29
rect -1356 8 -1354 29
rect -1348 8 -1346 29
rect -1340 8 -1338 29
rect -1332 8 -1330 29
rect -1300 26 -1298 28
rect -1300 13 -1298 23
rect -1266 25 -1264 32
rect -1258 25 -1256 32
rect -1250 25 -1248 32
rect -1242 25 -1240 32
rect -1234 25 -1232 32
rect -1181 25 -1179 32
rect -1173 25 -1171 32
rect -1165 25 -1163 32
rect -1157 25 -1155 32
rect -1149 25 -1147 32
rect -1141 25 -1139 32
rect -1133 25 -1131 32
rect -748 33 -746 40
rect -740 33 -738 40
rect -732 33 -730 40
rect -724 33 -722 40
rect -716 33 -714 40
rect -663 33 -661 40
rect -655 33 -653 40
rect -647 33 -645 40
rect -639 33 -637 40
rect -631 33 -629 40
rect -623 33 -621 40
rect -615 33 -613 40
rect -1642 -28 -1640 -26
rect -1642 -41 -1640 -31
rect -1465 -34 -1463 5
rect -1457 -4 -1455 5
rect -1449 -4 -1447 5
rect -1441 -4 -1439 5
rect -1433 -34 -1431 5
rect -1380 -4 -1378 5
rect -1372 -4 -1370 5
rect -1364 -4 -1362 5
rect -1356 -10 -1354 5
rect -1348 -4 -1346 5
rect -1340 -4 -1338 5
rect -1332 -4 -1330 5
rect -1300 2 -1298 10
rect -1266 1 -1264 22
rect -1258 1 -1256 22
rect -1250 1 -1248 22
rect -1242 1 -1240 22
rect -1234 1 -1232 22
rect -1181 1 -1179 22
rect -1173 1 -1171 22
rect -1165 1 -1163 22
rect -1157 1 -1155 22
rect -1149 1 -1147 22
rect -1141 1 -1139 22
rect -1133 1 -1131 22
rect -1101 19 -1099 21
rect -1063 19 -1061 26
rect -1055 19 -1053 26
rect -1047 19 -1045 26
rect -1039 19 -1037 26
rect -1031 19 -1029 26
rect -978 19 -976 26
rect -970 19 -968 26
rect -962 19 -960 26
rect -954 19 -952 26
rect -946 19 -944 26
rect -938 19 -936 26
rect -930 19 -928 26
rect -1101 6 -1099 16
rect -1388 -24 -1386 -22
rect -1388 -37 -1386 -27
rect -1266 -30 -1264 -2
rect -1258 -11 -1256 -2
rect -1250 -11 -1248 -2
rect -1242 -11 -1240 -2
rect -1234 -30 -1232 -2
rect -1181 -11 -1179 -2
rect -1173 -11 -1171 -2
rect -1165 -11 -1163 -2
rect -1157 -17 -1155 -2
rect -1149 -11 -1147 -2
rect -1141 -11 -1139 -2
rect -1133 -11 -1131 -2
rect -1101 -5 -1099 3
rect -1063 -5 -1061 16
rect -1055 -5 -1053 16
rect -1047 -5 -1045 16
rect -1039 -5 -1037 16
rect -1031 -5 -1029 16
rect -978 -5 -976 16
rect -970 -5 -968 16
rect -962 -5 -960 16
rect -954 -5 -952 16
rect -946 -5 -944 16
rect -938 -5 -936 16
rect -930 -5 -928 16
rect -898 13 -896 15
rect -898 0 -896 10
rect -748 9 -746 30
rect -740 9 -738 30
rect -732 9 -730 30
rect -724 9 -722 30
rect -716 9 -714 30
rect -663 9 -661 30
rect -655 9 -653 30
rect -647 9 -645 30
rect -639 9 -637 30
rect -631 9 -629 30
rect -623 9 -621 30
rect -615 9 -613 30
rect -583 27 -581 29
rect -583 14 -581 24
rect -495 24 -493 31
rect -487 24 -485 31
rect -479 24 -477 31
rect -471 24 -469 31
rect -463 24 -461 31
rect -410 24 -408 31
rect -402 24 -400 31
rect -394 24 -392 31
rect -386 24 -384 31
rect -378 24 -376 31
rect -370 24 -368 31
rect -362 24 -360 31
rect -1189 -31 -1187 -29
rect -1642 -52 -1640 -44
rect -1388 -48 -1386 -40
rect -1189 -44 -1187 -34
rect -1063 -37 -1061 -8
rect -1055 -17 -1053 -8
rect -1047 -17 -1045 -8
rect -1039 -17 -1037 -8
rect -1031 -37 -1029 -8
rect -978 -17 -976 -8
rect -970 -17 -968 -8
rect -962 -17 -960 -8
rect -954 -23 -952 -8
rect -946 -17 -944 -8
rect -938 -17 -936 -8
rect -930 -17 -928 -8
rect -898 -11 -896 -3
rect -986 -37 -984 -35
rect -1189 -55 -1187 -47
rect -986 -50 -984 -40
rect -748 -43 -746 6
rect -740 -3 -738 6
rect -732 -3 -730 6
rect -724 -3 -722 6
rect -716 -43 -714 6
rect -663 -3 -661 6
rect -655 -3 -653 6
rect -647 -3 -645 6
rect -639 -9 -637 6
rect -631 -3 -629 6
rect -623 -3 -621 6
rect -615 -3 -613 6
rect -583 3 -581 11
rect -495 0 -493 21
rect -487 0 -485 21
rect -479 0 -477 21
rect -471 0 -469 21
rect -463 0 -461 21
rect -410 0 -408 21
rect -402 0 -400 21
rect -394 0 -392 21
rect -386 0 -384 21
rect -378 0 -376 21
rect -370 0 -368 21
rect -362 0 -360 21
rect -330 18 -328 20
rect -252 18 -250 25
rect -244 18 -242 25
rect -236 18 -234 25
rect -228 18 -226 25
rect -220 18 -218 25
rect -167 18 -165 25
rect -159 18 -157 25
rect -151 18 -149 25
rect -143 18 -141 25
rect -135 18 -133 25
rect -127 18 -125 25
rect -119 18 -117 25
rect -330 5 -328 15
rect -671 -23 -669 -21
rect -671 -36 -669 -26
rect -495 -29 -493 -3
rect -487 -12 -485 -3
rect -479 -12 -477 -3
rect -471 -12 -469 -3
rect -463 -29 -461 -3
rect -410 -12 -408 -3
rect -402 -12 -400 -3
rect -394 -12 -392 -3
rect -386 -18 -384 -3
rect -378 -12 -376 -3
rect -370 -12 -368 -3
rect -362 -12 -360 -3
rect -330 -6 -328 2
rect -252 -6 -250 15
rect -244 -6 -242 15
rect -236 -6 -234 15
rect -228 -6 -226 15
rect -220 -6 -218 15
rect -167 -6 -165 15
rect -159 -6 -157 15
rect -151 -6 -149 15
rect -143 -6 -141 15
rect -135 -6 -133 15
rect -127 -6 -125 15
rect -119 -6 -117 15
rect -87 12 -85 14
rect -6 14 -4 21
rect 2 14 4 21
rect 10 14 12 21
rect 18 14 20 21
rect 26 14 28 21
rect 79 14 81 21
rect 87 14 89 21
rect 95 14 97 21
rect 103 14 105 21
rect 111 14 113 21
rect 119 14 121 21
rect 127 14 129 21
rect -87 -1 -85 9
rect -418 -32 -416 -30
rect -671 -47 -669 -39
rect -418 -45 -416 -35
rect -252 -38 -250 -9
rect -244 -18 -242 -9
rect -236 -18 -234 -9
rect -228 -18 -226 -9
rect -220 -38 -218 -9
rect -167 -18 -165 -9
rect -159 -18 -157 -9
rect -151 -18 -149 -9
rect -143 -24 -141 -9
rect -135 -18 -133 -9
rect -127 -18 -125 -9
rect -119 -18 -117 -9
rect -87 -12 -85 -4
rect -6 -10 -4 11
rect 2 -10 4 11
rect 10 -10 12 11
rect 18 -10 20 11
rect 26 -10 28 11
rect 79 -10 81 11
rect 87 -10 89 11
rect 95 -10 97 11
rect 103 -10 105 11
rect 111 -10 113 11
rect 119 -10 121 11
rect 127 -10 129 11
rect 159 8 161 10
rect 159 -5 161 5
rect -175 -38 -173 -36
rect -986 -61 -984 -53
rect -418 -56 -416 -48
rect -175 -51 -173 -41
rect -6 -44 -4 -13
rect 2 -22 4 -13
rect 10 -22 12 -13
rect 18 -22 20 -13
rect 26 -44 28 -13
rect 79 -22 81 -13
rect 87 -22 89 -13
rect 95 -22 97 -13
rect 103 -28 105 -13
rect 111 -22 113 -13
rect 119 -22 121 -13
rect 127 -22 129 -13
rect 159 -16 161 -8
rect 71 -42 73 -40
rect -175 -62 -173 -54
rect 71 -55 73 -45
rect 71 -66 73 -58
<< ndiffusion >>
rect -1555 6 -1554 9
rect -1552 6 -1551 9
rect -1720 1 -1719 4
rect -1717 1 -1711 4
rect -1709 1 -1708 4
rect -1704 1 -1703 4
rect -1701 1 -1700 4
rect -1696 1 -1695 4
rect -1693 1 -1692 4
rect -1688 1 -1687 4
rect -1685 1 -1684 4
rect -1635 1 -1634 4
rect -1632 1 -1631 4
rect -1627 1 -1626 4
rect -1624 1 -1623 4
rect -1619 1 -1618 4
rect -1616 1 -1615 4
rect -1611 1 -1610 4
rect -1608 1 -1607 4
rect -1603 1 -1602 4
rect -1600 1 -1594 4
rect -1592 1 -1586 4
rect -1584 1 -1583 4
rect -1301 10 -1300 13
rect -1298 10 -1297 13
rect -1466 5 -1465 8
rect -1463 5 -1457 8
rect -1455 5 -1454 8
rect -1450 5 -1449 8
rect -1447 5 -1446 8
rect -1442 5 -1441 8
rect -1439 5 -1438 8
rect -1434 5 -1433 8
rect -1431 5 -1430 8
rect -1381 5 -1380 8
rect -1378 5 -1377 8
rect -1373 5 -1372 8
rect -1370 5 -1369 8
rect -1365 5 -1364 8
rect -1362 5 -1361 8
rect -1357 5 -1356 8
rect -1354 5 -1353 8
rect -1349 5 -1348 8
rect -1346 5 -1340 8
rect -1338 5 -1332 8
rect -1330 5 -1329 8
rect -1102 3 -1101 6
rect -1099 3 -1098 6
rect -1267 -2 -1266 1
rect -1264 -2 -1258 1
rect -1256 -2 -1255 1
rect -1251 -2 -1250 1
rect -1248 -2 -1247 1
rect -1243 -2 -1242 1
rect -1240 -2 -1239 1
rect -1235 -2 -1234 1
rect -1232 -2 -1231 1
rect -1182 -2 -1181 1
rect -1179 -2 -1178 1
rect -1174 -2 -1173 1
rect -1171 -2 -1170 1
rect -1166 -2 -1165 1
rect -1163 -2 -1162 1
rect -1158 -2 -1157 1
rect -1155 -2 -1154 1
rect -1150 -2 -1149 1
rect -1147 -2 -1141 1
rect -1139 -2 -1133 1
rect -1131 -2 -1130 1
rect -584 11 -583 14
rect -581 11 -580 14
rect -749 6 -748 9
rect -746 6 -740 9
rect -738 6 -737 9
rect -899 -3 -898 0
rect -896 -3 -895 0
rect -1064 -8 -1063 -5
rect -1061 -8 -1055 -5
rect -1053 -8 -1052 -5
rect -1389 -40 -1388 -37
rect -1386 -40 -1385 -37
rect -1643 -44 -1642 -41
rect -1640 -44 -1639 -41
rect -1048 -8 -1047 -5
rect -1045 -8 -1044 -5
rect -1040 -8 -1039 -5
rect -1037 -8 -1036 -5
rect -1032 -8 -1031 -5
rect -1029 -8 -1028 -5
rect -979 -8 -978 -5
rect -976 -8 -975 -5
rect -971 -8 -970 -5
rect -968 -8 -967 -5
rect -963 -8 -962 -5
rect -960 -8 -959 -5
rect -955 -8 -954 -5
rect -952 -8 -951 -5
rect -947 -8 -946 -5
rect -944 -8 -938 -5
rect -936 -8 -930 -5
rect -928 -8 -927 -5
rect -1190 -47 -1189 -44
rect -1187 -47 -1186 -44
rect -733 6 -732 9
rect -730 6 -729 9
rect -725 6 -724 9
rect -722 6 -721 9
rect -717 6 -716 9
rect -714 6 -713 9
rect -664 6 -663 9
rect -661 6 -660 9
rect -656 6 -655 9
rect -653 6 -652 9
rect -648 6 -647 9
rect -645 6 -644 9
rect -640 6 -639 9
rect -637 6 -636 9
rect -632 6 -631 9
rect -629 6 -623 9
rect -621 6 -615 9
rect -613 6 -612 9
rect -331 2 -330 5
rect -328 2 -327 5
rect -496 -3 -495 0
rect -493 -3 -487 0
rect -485 -3 -484 0
rect -480 -3 -479 0
rect -477 -3 -476 0
rect -472 -3 -471 0
rect -469 -3 -468 0
rect -464 -3 -463 0
rect -461 -3 -460 0
rect -411 -3 -410 0
rect -408 -3 -407 0
rect -403 -3 -402 0
rect -400 -3 -399 0
rect -395 -3 -394 0
rect -392 -3 -391 0
rect -387 -3 -386 0
rect -384 -3 -383 0
rect -379 -3 -378 0
rect -376 -3 -370 0
rect -368 -3 -362 0
rect -360 -3 -359 0
rect -88 -4 -87 -1
rect -85 -4 -84 -1
rect -253 -9 -252 -6
rect -250 -9 -244 -6
rect -242 -9 -241 -6
rect -672 -39 -671 -36
rect -669 -39 -668 -36
rect -237 -9 -236 -6
rect -234 -9 -233 -6
rect -229 -9 -228 -6
rect -226 -9 -225 -6
rect -221 -9 -220 -6
rect -218 -9 -217 -6
rect -168 -9 -167 -6
rect -165 -9 -164 -6
rect -160 -9 -159 -6
rect -157 -9 -156 -6
rect -152 -9 -151 -6
rect -149 -9 -148 -6
rect -144 -9 -143 -6
rect -141 -9 -140 -6
rect -136 -9 -135 -6
rect -133 -9 -127 -6
rect -125 -9 -119 -6
rect -117 -9 -116 -6
rect 158 -8 159 -5
rect 161 -8 162 -5
rect -7 -13 -6 -10
rect -4 -13 2 -10
rect 4 -13 5 -10
rect -419 -48 -418 -45
rect -416 -48 -415 -45
rect -987 -53 -986 -50
rect -984 -53 -983 -50
rect 9 -13 10 -10
rect 12 -13 13 -10
rect 17 -13 18 -10
rect 20 -13 21 -10
rect 25 -13 26 -10
rect 28 -13 29 -10
rect 78 -13 79 -10
rect 81 -13 82 -10
rect 86 -13 87 -10
rect 89 -13 90 -10
rect 94 -13 95 -10
rect 97 -13 98 -10
rect 102 -13 103 -10
rect 105 -13 106 -10
rect 110 -13 111 -10
rect 113 -13 119 -10
rect 121 -13 127 -10
rect 129 -13 130 -10
rect -176 -54 -175 -51
rect -173 -54 -172 -51
rect 70 -58 71 -55
rect 73 -58 74 -55
<< pdiffusion >>
rect -1720 25 -1719 28
rect -1717 25 -1716 28
rect -1712 25 -1711 28
rect -1709 25 -1708 28
rect -1704 25 -1703 28
rect -1701 25 -1700 28
rect -1696 25 -1695 28
rect -1693 25 -1687 28
rect -1685 25 -1684 28
rect -1635 25 -1634 28
rect -1632 25 -1626 28
rect -1624 25 -1618 28
rect -1616 25 -1615 28
rect -1611 25 -1610 28
rect -1608 25 -1607 28
rect -1603 25 -1602 28
rect -1600 25 -1599 28
rect -1595 25 -1594 28
rect -1592 25 -1591 28
rect -1587 25 -1586 28
rect -1584 25 -1583 28
rect -1466 29 -1465 32
rect -1463 29 -1462 32
rect -1458 29 -1457 32
rect -1455 29 -1454 32
rect -1450 29 -1449 32
rect -1447 29 -1446 32
rect -1442 29 -1441 32
rect -1439 29 -1433 32
rect -1431 29 -1430 32
rect -1381 29 -1380 32
rect -1378 29 -1372 32
rect -1370 29 -1364 32
rect -1362 29 -1361 32
rect -1357 29 -1356 32
rect -1354 29 -1353 32
rect -1349 29 -1348 32
rect -1346 29 -1345 32
rect -1341 29 -1340 32
rect -1338 29 -1337 32
rect -1333 29 -1332 32
rect -1330 29 -1329 32
rect -1555 19 -1554 22
rect -1552 19 -1551 22
rect -1301 23 -1300 26
rect -1298 23 -1297 26
rect -1267 22 -1266 25
rect -1264 22 -1263 25
rect -1259 22 -1258 25
rect -1256 22 -1255 25
rect -1251 22 -1250 25
rect -1248 22 -1247 25
rect -1243 22 -1242 25
rect -1240 22 -1234 25
rect -1232 22 -1231 25
rect -1182 22 -1181 25
rect -1179 22 -1173 25
rect -1171 22 -1165 25
rect -1163 22 -1162 25
rect -1158 22 -1157 25
rect -1155 22 -1154 25
rect -1150 22 -1149 25
rect -1147 22 -1146 25
rect -1142 22 -1141 25
rect -1139 22 -1138 25
rect -749 30 -748 33
rect -746 30 -745 33
rect -741 30 -740 33
rect -738 30 -737 33
rect -733 30 -732 33
rect -730 30 -729 33
rect -725 30 -724 33
rect -722 30 -716 33
rect -714 30 -713 33
rect -664 30 -663 33
rect -661 30 -655 33
rect -653 30 -647 33
rect -645 30 -644 33
rect -640 30 -639 33
rect -637 30 -636 33
rect -632 30 -631 33
rect -629 30 -628 33
rect -624 30 -623 33
rect -621 30 -620 33
rect -616 30 -615 33
rect -613 30 -612 33
rect -1134 22 -1133 25
rect -1131 22 -1130 25
rect -1643 -31 -1642 -28
rect -1640 -31 -1639 -28
rect -1102 16 -1101 19
rect -1099 16 -1098 19
rect -1064 16 -1063 19
rect -1061 16 -1060 19
rect -1056 16 -1055 19
rect -1053 16 -1052 19
rect -1048 16 -1047 19
rect -1045 16 -1044 19
rect -1040 16 -1039 19
rect -1037 16 -1031 19
rect -1029 16 -1028 19
rect -979 16 -978 19
rect -976 16 -970 19
rect -968 16 -962 19
rect -960 16 -959 19
rect -955 16 -954 19
rect -952 16 -951 19
rect -947 16 -946 19
rect -944 16 -943 19
rect -939 16 -938 19
rect -936 16 -935 19
rect -931 16 -930 19
rect -928 16 -927 19
rect -1389 -27 -1388 -24
rect -1386 -27 -1385 -24
rect -899 10 -898 13
rect -896 10 -895 13
rect -584 24 -583 27
rect -581 24 -580 27
rect -496 21 -495 24
rect -493 21 -492 24
rect -488 21 -487 24
rect -485 21 -484 24
rect -480 21 -479 24
rect -477 21 -476 24
rect -472 21 -471 24
rect -469 21 -463 24
rect -461 21 -460 24
rect -411 21 -410 24
rect -408 21 -402 24
rect -400 21 -394 24
rect -392 21 -391 24
rect -387 21 -386 24
rect -384 21 -383 24
rect -379 21 -378 24
rect -376 21 -375 24
rect -371 21 -370 24
rect -368 21 -367 24
rect -363 21 -362 24
rect -360 21 -359 24
rect -1190 -34 -1189 -31
rect -1187 -34 -1186 -31
rect -987 -40 -986 -37
rect -984 -40 -983 -37
rect -331 15 -330 18
rect -328 15 -327 18
rect -253 15 -252 18
rect -250 15 -249 18
rect -245 15 -244 18
rect -242 15 -241 18
rect -237 15 -236 18
rect -234 15 -233 18
rect -229 15 -228 18
rect -226 15 -220 18
rect -218 15 -217 18
rect -168 15 -167 18
rect -165 15 -159 18
rect -157 15 -151 18
rect -149 15 -148 18
rect -144 15 -143 18
rect -141 15 -140 18
rect -136 15 -135 18
rect -133 15 -132 18
rect -128 15 -127 18
rect -125 15 -124 18
rect -120 15 -119 18
rect -117 15 -116 18
rect -672 -26 -671 -23
rect -669 -26 -668 -23
rect -88 9 -87 12
rect -85 9 -84 12
rect -7 11 -6 14
rect -4 11 -3 14
rect 1 11 2 14
rect 4 11 5 14
rect 9 11 10 14
rect 12 11 13 14
rect 17 11 18 14
rect 20 11 26 14
rect 28 11 29 14
rect 78 11 79 14
rect 81 11 87 14
rect 89 11 95 14
rect 97 11 98 14
rect 102 11 103 14
rect 105 11 106 14
rect 110 11 111 14
rect 113 11 114 14
rect 118 11 119 14
rect 121 11 122 14
rect 126 11 127 14
rect 129 11 130 14
rect -419 -35 -418 -32
rect -416 -35 -415 -32
rect 158 5 159 8
rect 161 5 162 8
rect -176 -41 -175 -38
rect -173 -41 -172 -38
rect 70 -45 71 -42
rect 73 -45 74 -42
<< metal1 >>
rect -1472 42 -1446 45
rect -1442 42 -1424 45
rect -1387 42 -1361 45
rect -1726 38 -1700 41
rect -1696 38 -1678 41
rect -1641 38 -1615 41
rect -1724 32 -1705 35
rect -1724 29 -1721 32
rect -1708 29 -1705 32
rect -1699 29 -1696 38
rect -1611 38 -1577 41
rect -1614 29 -1611 37
rect -1470 36 -1451 39
rect -1716 16 -1713 25
rect -1708 22 -1705 25
rect -1683 22 -1680 25
rect -1708 19 -1680 22
rect -1607 32 -1587 35
rect -1607 29 -1604 32
rect -1590 29 -1587 32
rect -1470 33 -1467 36
rect -1454 33 -1451 36
rect -1445 33 -1442 42
rect -1357 42 -1323 45
rect -755 43 -729 46
rect -725 43 -707 46
rect -670 43 -644 46
rect -1360 33 -1357 41
rect -1639 22 -1636 25
rect -1606 22 -1603 25
rect -1639 19 -1603 22
rect -1598 16 -1595 25
rect -1582 16 -1579 25
rect -1555 27 -1547 30
rect -1559 23 -1556 27
rect -1462 20 -1459 29
rect -1454 26 -1451 29
rect -1429 26 -1426 29
rect -1454 23 -1426 26
rect -1353 36 -1333 39
rect -1353 33 -1350 36
rect -1336 33 -1333 36
rect -1273 35 -1247 38
rect -1243 35 -1225 38
rect -1188 35 -1162 38
rect -1385 26 -1382 29
rect -1352 26 -1349 29
rect -1385 23 -1349 26
rect -1344 20 -1341 29
rect -1328 20 -1325 29
rect -1301 31 -1293 34
rect -1305 27 -1302 31
rect -1271 29 -1252 32
rect -1296 20 -1293 23
rect -1271 26 -1268 29
rect -1255 26 -1252 29
rect -1246 26 -1243 35
rect -1158 35 -1124 38
rect -753 37 -734 40
rect -1161 26 -1158 34
rect -753 34 -750 37
rect -737 34 -734 37
rect -728 34 -725 43
rect -640 43 -606 46
rect -643 34 -640 42
rect -1550 16 -1547 19
rect -1472 17 -1405 20
rect -1387 17 -1304 20
rect -1726 13 -1659 16
rect -1641 13 -1558 16
rect -1708 4 -1705 13
rect -1700 7 -1680 10
rect -1700 4 -1697 7
rect -1683 4 -1680 7
rect -1724 -4 -1721 0
rect -1691 -4 -1688 0
rect -1726 -8 -1725 -5
rect -1721 -8 -1692 -5
rect -1688 -8 -1678 -5
rect -1662 -11 -1659 13
rect -1631 7 -1611 10
rect -1631 4 -1628 7
rect -1614 4 -1611 7
rect -1607 4 -1604 13
rect -1550 13 -1538 16
rect -1550 9 -1547 13
rect -1454 8 -1451 17
rect -1446 11 -1426 14
rect -1446 8 -1443 11
rect -1429 8 -1426 11
rect -1639 -4 -1636 0
rect -1622 -4 -1619 0
rect -1641 -8 -1640 -5
rect -1636 -8 -1623 -5
rect -1582 -4 -1579 0
rect -1559 1 -1556 5
rect -1555 -2 -1547 1
rect -1470 0 -1467 4
rect -1437 0 -1434 4
rect -1472 -4 -1471 -1
rect -1467 -4 -1438 -1
rect -1434 -4 -1424 -1
rect -1619 -8 -1582 -5
rect -1578 -8 -1577 -5
rect -1408 -7 -1405 17
rect -1377 11 -1357 14
rect -1377 8 -1374 11
rect -1360 8 -1357 11
rect -1353 8 -1350 17
rect -1296 17 -1284 20
rect -1296 13 -1293 17
rect -1263 13 -1260 22
rect -1255 19 -1252 22
rect -1230 19 -1227 22
rect -1255 16 -1227 19
rect -1154 29 -1134 32
rect -1070 29 -1044 32
rect -1040 29 -1022 32
rect -985 29 -959 32
rect -1154 26 -1151 29
rect -1137 26 -1134 29
rect -1186 19 -1183 22
rect -1153 19 -1150 22
rect -1186 16 -1150 19
rect -1145 13 -1142 22
rect -1129 13 -1126 22
rect -1102 24 -1094 27
rect -1106 20 -1103 24
rect -1068 23 -1049 26
rect -1068 20 -1065 23
rect -1052 20 -1049 23
rect -1043 20 -1040 29
rect -955 29 -921 32
rect -958 20 -955 28
rect -1097 13 -1094 16
rect -1273 10 -1206 13
rect -1188 10 -1105 13
rect -1385 0 -1382 4
rect -1368 0 -1365 4
rect -1387 -4 -1386 -1
rect -1382 -4 -1369 -1
rect -1328 0 -1325 4
rect -1305 5 -1302 9
rect -1301 2 -1293 5
rect -1255 1 -1252 10
rect -1247 4 -1227 7
rect -1247 1 -1244 4
rect -1230 1 -1227 4
rect -1365 -4 -1328 -1
rect -1324 -4 -1323 -1
rect -1271 -7 -1268 -3
rect -1238 -7 -1235 -3
rect -1408 -10 -1360 -7
rect -1662 -14 -1614 -11
rect -1662 -35 -1659 -14
rect -1643 -23 -1635 -20
rect -1647 -27 -1644 -23
rect -1638 -34 -1635 -31
rect -1408 -31 -1405 -10
rect -1273 -11 -1272 -8
rect -1268 -11 -1239 -8
rect -1235 -11 -1225 -8
rect -1209 -14 -1206 10
rect -1178 4 -1158 7
rect -1178 1 -1175 4
rect -1161 1 -1158 4
rect -1154 1 -1151 10
rect -1097 10 -1085 13
rect -1097 6 -1094 10
rect -1060 7 -1057 16
rect -1052 13 -1049 16
rect -1027 13 -1024 16
rect -1052 10 -1024 13
rect -951 23 -931 26
rect -951 20 -948 23
rect -934 20 -931 23
rect -983 13 -980 16
rect -950 13 -947 16
rect -983 10 -947 13
rect -942 7 -939 16
rect -926 7 -923 16
rect -745 21 -742 30
rect -737 27 -734 30
rect -712 27 -709 30
rect -737 24 -709 27
rect -636 37 -616 40
rect -636 34 -633 37
rect -619 34 -616 37
rect -668 27 -665 30
rect -635 27 -632 30
rect -668 24 -632 27
rect -627 21 -624 30
rect -611 21 -608 30
rect -584 32 -576 35
rect -502 34 -476 37
rect -472 34 -454 37
rect -417 34 -391 37
rect -588 28 -585 32
rect -500 28 -481 31
rect -579 21 -576 24
rect -500 25 -497 28
rect -484 25 -481 28
rect -475 25 -472 34
rect -387 34 -353 37
rect -390 25 -387 33
rect -899 18 -891 21
rect -755 18 -688 21
rect -670 18 -587 21
rect -903 14 -900 18
rect -894 7 -891 10
rect -737 9 -734 18
rect -729 12 -709 15
rect -729 9 -726 12
rect -712 9 -709 12
rect -1070 4 -1003 7
rect -985 4 -902 7
rect -1186 -7 -1183 -3
rect -1169 -7 -1166 -3
rect -1188 -11 -1187 -8
rect -1183 -11 -1170 -8
rect -1129 -7 -1126 -3
rect -1106 -2 -1103 2
rect -1102 -5 -1094 -2
rect -1052 -5 -1049 4
rect -1044 -2 -1024 1
rect -1044 -5 -1041 -2
rect -1027 -5 -1024 -2
rect -1166 -11 -1129 -8
rect -1125 -11 -1124 -8
rect -1068 -13 -1065 -9
rect -1035 -13 -1032 -9
rect -1389 -19 -1381 -16
rect -1209 -17 -1161 -14
rect -1393 -23 -1390 -19
rect -1384 -30 -1381 -27
rect -1408 -34 -1392 -31
rect -1384 -33 -1267 -30
rect -1662 -38 -1646 -35
rect -1638 -37 -1466 -34
rect -1638 -41 -1635 -37
rect -1462 -37 -1434 -34
rect -1384 -37 -1381 -33
rect -1263 -33 -1235 -30
rect -1209 -38 -1206 -17
rect -1070 -17 -1069 -14
rect -1065 -17 -1036 -14
rect -1032 -17 -1022 -14
rect -1006 -20 -1003 4
rect -975 -2 -955 1
rect -975 -5 -972 -2
rect -958 -5 -955 -2
rect -951 -5 -948 4
rect -894 4 -882 7
rect -894 0 -891 4
rect -753 1 -750 5
rect -720 1 -717 5
rect -755 -3 -754 0
rect -750 -3 -721 0
rect -717 -3 -707 0
rect -983 -13 -980 -9
rect -966 -13 -963 -9
rect -985 -17 -984 -14
rect -980 -17 -967 -14
rect -926 -13 -923 -9
rect -903 -8 -900 -4
rect -691 -6 -688 18
rect -660 12 -640 15
rect -660 9 -657 12
rect -643 9 -640 12
rect -636 9 -633 18
rect -579 18 -567 21
rect -579 14 -576 18
rect -492 12 -489 21
rect -484 18 -481 21
rect -459 18 -456 21
rect -484 15 -456 18
rect -383 28 -363 31
rect -259 28 -233 31
rect -229 28 -211 31
rect -174 28 -148 31
rect -383 25 -380 28
rect -366 25 -363 28
rect -415 18 -412 21
rect -382 18 -379 21
rect -415 15 -379 18
rect -374 12 -371 21
rect -358 12 -355 21
rect -331 23 -323 26
rect -335 19 -332 23
rect -257 22 -238 25
rect -257 19 -254 22
rect -241 19 -238 22
rect -232 19 -229 28
rect -144 28 -110 31
rect -147 19 -144 27
rect -326 12 -323 15
rect -668 1 -665 5
rect -651 1 -648 5
rect -670 -3 -669 0
rect -665 -3 -652 0
rect -611 1 -608 5
rect -588 6 -585 10
rect -502 9 -435 12
rect -417 9 -334 12
rect -584 3 -576 6
rect -648 -3 -611 0
rect -484 0 -481 9
rect -476 3 -456 6
rect -476 0 -473 3
rect -459 0 -456 3
rect -607 -3 -606 0
rect -899 -11 -891 -8
rect -691 -9 -643 -6
rect -963 -17 -926 -14
rect -922 -17 -921 -14
rect -1006 -23 -958 -20
rect -1190 -26 -1182 -23
rect -1194 -30 -1191 -26
rect -1185 -37 -1182 -34
rect -1209 -41 -1193 -38
rect -1185 -40 -1064 -37
rect -1393 -45 -1390 -41
rect -1185 -44 -1182 -40
rect -1060 -40 -1032 -37
rect -1028 -40 -1027 -37
rect -1647 -49 -1644 -45
rect -1389 -48 -1381 -45
rect -1006 -44 -1003 -23
rect -987 -32 -979 -29
rect -691 -30 -688 -9
rect -500 -8 -497 -4
rect -467 -8 -464 -4
rect -502 -12 -501 -9
rect -497 -12 -468 -9
rect -464 -12 -454 -9
rect -438 -15 -435 9
rect -407 3 -387 6
rect -407 0 -404 3
rect -390 0 -387 3
rect -383 0 -380 9
rect -326 9 -314 12
rect -326 5 -323 9
rect -249 6 -246 15
rect -241 12 -238 15
rect -216 12 -213 15
rect -241 9 -213 12
rect -140 22 -120 25
rect -13 24 13 27
rect 17 24 35 27
rect 72 24 98 27
rect -140 19 -137 22
rect -123 19 -120 22
rect -172 12 -169 15
rect -139 12 -136 15
rect -172 9 -136 12
rect -131 6 -128 15
rect -115 6 -112 15
rect -88 17 -80 20
rect -11 18 8 21
rect -92 13 -89 17
rect -11 15 -8 18
rect 5 15 8 18
rect 14 15 17 24
rect 102 24 136 27
rect 99 15 102 23
rect -83 6 -80 9
rect -259 3 -192 6
rect -174 3 -91 6
rect -415 -8 -412 -4
rect -398 -8 -395 -4
rect -417 -12 -416 -9
rect -412 -12 -399 -9
rect -358 -8 -355 -4
rect -335 -3 -332 1
rect -331 -6 -323 -3
rect -241 -6 -238 3
rect -233 -3 -213 0
rect -233 -6 -230 -3
rect -216 -6 -213 -3
rect -395 -12 -358 -9
rect -354 -12 -353 -9
rect -257 -14 -254 -10
rect -224 -14 -221 -10
rect -672 -18 -664 -15
rect -438 -18 -390 -15
rect -676 -22 -673 -18
rect -667 -29 -664 -26
rect -991 -36 -988 -32
rect -691 -33 -675 -30
rect -667 -32 -496 -29
rect -667 -36 -664 -32
rect -492 -32 -464 -29
rect -982 -43 -979 -40
rect -438 -39 -435 -18
rect -259 -18 -258 -15
rect -254 -18 -225 -15
rect -221 -18 -211 -15
rect -195 -21 -192 3
rect -164 -3 -144 0
rect -164 -6 -161 -3
rect -147 -6 -144 -3
rect -140 -6 -137 3
rect -83 3 -71 6
rect -83 -1 -80 3
rect -3 2 0 11
rect 5 8 8 11
rect 30 8 33 11
rect 5 5 33 8
rect 106 18 126 21
rect 106 15 109 18
rect 123 15 126 18
rect 74 8 77 11
rect 107 8 110 11
rect 74 5 110 8
rect 115 2 118 11
rect 131 2 134 11
rect 158 13 166 16
rect 154 9 157 13
rect 163 2 166 5
rect -13 -1 54 2
rect 72 -1 155 2
rect -172 -14 -169 -10
rect -155 -14 -152 -10
rect -174 -18 -173 -15
rect -169 -18 -156 -15
rect -115 -14 -112 -10
rect -92 -9 -89 -5
rect -88 -12 -80 -9
rect 5 -10 8 -1
rect 13 -7 33 -4
rect 13 -10 16 -7
rect 30 -10 33 -7
rect -152 -18 -115 -15
rect -111 -18 -110 -15
rect -11 -18 -8 -14
rect 22 -18 25 -14
rect -195 -24 -147 -21
rect -419 -27 -411 -24
rect -423 -31 -420 -27
rect -414 -38 -411 -35
rect -1006 -47 -990 -44
rect -982 -46 -749 -43
rect -1643 -52 -1635 -49
rect -1194 -52 -1191 -48
rect -982 -50 -979 -46
rect -745 -46 -717 -43
rect -676 -44 -673 -40
rect -438 -42 -422 -39
rect -414 -41 -253 -38
rect -672 -47 -664 -44
rect -414 -45 -411 -41
rect -249 -41 -221 -38
rect -1190 -55 -1182 -52
rect -195 -45 -192 -24
rect -13 -22 -12 -19
rect -8 -22 21 -19
rect 25 -22 35 -19
rect 51 -25 54 -1
rect 82 -7 102 -4
rect 82 -10 85 -7
rect 99 -10 102 -7
rect 106 -10 109 -1
rect 163 -1 175 2
rect 163 -5 166 -1
rect 74 -18 77 -14
rect 91 -18 94 -14
rect 72 -22 73 -19
rect 77 -22 90 -19
rect 131 -18 134 -14
rect 154 -13 157 -9
rect 158 -16 166 -13
rect 94 -22 131 -19
rect 135 -22 136 -19
rect 51 -28 99 -25
rect -176 -33 -168 -30
rect -180 -37 -177 -33
rect -171 -44 -168 -41
rect -195 -48 -179 -45
rect -171 -47 -7 -44
rect -423 -53 -420 -49
rect -171 -51 -168 -47
rect -3 -47 25 -44
rect -991 -58 -988 -54
rect -419 -56 -411 -53
rect 51 -49 54 -28
rect 70 -37 78 -34
rect 66 -41 69 -37
rect 75 -48 78 -45
rect 51 -52 67 -49
rect 75 -51 86 -48
rect 75 -55 78 -51
rect -987 -61 -979 -58
rect -180 -59 -177 -55
rect -176 -62 -168 -59
rect 66 -63 69 -59
rect 70 -66 78 -63
<< ntransistor >>
rect -1554 6 -1552 9
rect -1719 1 -1717 4
rect -1711 1 -1709 4
rect -1703 1 -1701 4
rect -1695 1 -1693 4
rect -1687 1 -1685 4
rect -1634 1 -1632 4
rect -1626 1 -1624 4
rect -1618 1 -1616 4
rect -1610 1 -1608 4
rect -1602 1 -1600 4
rect -1594 1 -1592 4
rect -1586 1 -1584 4
rect -1300 10 -1298 13
rect -1465 5 -1463 8
rect -1457 5 -1455 8
rect -1449 5 -1447 8
rect -1441 5 -1439 8
rect -1433 5 -1431 8
rect -1380 5 -1378 8
rect -1372 5 -1370 8
rect -1364 5 -1362 8
rect -1356 5 -1354 8
rect -1348 5 -1346 8
rect -1340 5 -1338 8
rect -1332 5 -1330 8
rect -1101 3 -1099 6
rect -1266 -2 -1264 1
rect -1258 -2 -1256 1
rect -1250 -2 -1248 1
rect -1242 -2 -1240 1
rect -1234 -2 -1232 1
rect -1181 -2 -1179 1
rect -1173 -2 -1171 1
rect -1165 -2 -1163 1
rect -1157 -2 -1155 1
rect -1149 -2 -1147 1
rect -1141 -2 -1139 1
rect -1133 -2 -1131 1
rect -583 11 -581 14
rect -748 6 -746 9
rect -740 6 -738 9
rect -898 -3 -896 0
rect -1063 -8 -1061 -5
rect -1055 -8 -1053 -5
rect -1388 -40 -1386 -37
rect -1642 -44 -1640 -41
rect -1047 -8 -1045 -5
rect -1039 -8 -1037 -5
rect -1031 -8 -1029 -5
rect -978 -8 -976 -5
rect -970 -8 -968 -5
rect -962 -8 -960 -5
rect -954 -8 -952 -5
rect -946 -8 -944 -5
rect -938 -8 -936 -5
rect -930 -8 -928 -5
rect -1189 -47 -1187 -44
rect -732 6 -730 9
rect -724 6 -722 9
rect -716 6 -714 9
rect -663 6 -661 9
rect -655 6 -653 9
rect -647 6 -645 9
rect -639 6 -637 9
rect -631 6 -629 9
rect -623 6 -621 9
rect -615 6 -613 9
rect -330 2 -328 5
rect -495 -3 -493 0
rect -487 -3 -485 0
rect -479 -3 -477 0
rect -471 -3 -469 0
rect -463 -3 -461 0
rect -410 -3 -408 0
rect -402 -3 -400 0
rect -394 -3 -392 0
rect -386 -3 -384 0
rect -378 -3 -376 0
rect -370 -3 -368 0
rect -362 -3 -360 0
rect -87 -4 -85 -1
rect -252 -9 -250 -6
rect -244 -9 -242 -6
rect -671 -39 -669 -36
rect -236 -9 -234 -6
rect -228 -9 -226 -6
rect -220 -9 -218 -6
rect -167 -9 -165 -6
rect -159 -9 -157 -6
rect -151 -9 -149 -6
rect -143 -9 -141 -6
rect -135 -9 -133 -6
rect -127 -9 -125 -6
rect -119 -9 -117 -6
rect 159 -8 161 -5
rect -6 -13 -4 -10
rect 2 -13 4 -10
rect -418 -48 -416 -45
rect -986 -53 -984 -50
rect 10 -13 12 -10
rect 18 -13 20 -10
rect 26 -13 28 -10
rect 79 -13 81 -10
rect 87 -13 89 -10
rect 95 -13 97 -10
rect 103 -13 105 -10
rect 111 -13 113 -10
rect 119 -13 121 -10
rect 127 -13 129 -10
rect -175 -54 -173 -51
rect 71 -58 73 -55
<< ptransistor >>
rect -1719 25 -1717 28
rect -1711 25 -1709 28
rect -1703 25 -1701 28
rect -1695 25 -1693 28
rect -1687 25 -1685 28
rect -1634 25 -1632 28
rect -1626 25 -1624 28
rect -1618 25 -1616 28
rect -1610 25 -1608 28
rect -1602 25 -1600 28
rect -1594 25 -1592 28
rect -1586 25 -1584 28
rect -1465 29 -1463 32
rect -1457 29 -1455 32
rect -1449 29 -1447 32
rect -1441 29 -1439 32
rect -1433 29 -1431 32
rect -1380 29 -1378 32
rect -1372 29 -1370 32
rect -1364 29 -1362 32
rect -1356 29 -1354 32
rect -1348 29 -1346 32
rect -1340 29 -1338 32
rect -1332 29 -1330 32
rect -1554 19 -1552 22
rect -1300 23 -1298 26
rect -1266 22 -1264 25
rect -1258 22 -1256 25
rect -1250 22 -1248 25
rect -1242 22 -1240 25
rect -1234 22 -1232 25
rect -1181 22 -1179 25
rect -1173 22 -1171 25
rect -1165 22 -1163 25
rect -1157 22 -1155 25
rect -1149 22 -1147 25
rect -1141 22 -1139 25
rect -748 30 -746 33
rect -740 30 -738 33
rect -732 30 -730 33
rect -724 30 -722 33
rect -716 30 -714 33
rect -663 30 -661 33
rect -655 30 -653 33
rect -647 30 -645 33
rect -639 30 -637 33
rect -631 30 -629 33
rect -623 30 -621 33
rect -615 30 -613 33
rect -1133 22 -1131 25
rect -1642 -31 -1640 -28
rect -1101 16 -1099 19
rect -1063 16 -1061 19
rect -1055 16 -1053 19
rect -1047 16 -1045 19
rect -1039 16 -1037 19
rect -1031 16 -1029 19
rect -978 16 -976 19
rect -970 16 -968 19
rect -962 16 -960 19
rect -954 16 -952 19
rect -946 16 -944 19
rect -938 16 -936 19
rect -930 16 -928 19
rect -1388 -27 -1386 -24
rect -898 10 -896 13
rect -583 24 -581 27
rect -495 21 -493 24
rect -487 21 -485 24
rect -479 21 -477 24
rect -471 21 -469 24
rect -463 21 -461 24
rect -410 21 -408 24
rect -402 21 -400 24
rect -394 21 -392 24
rect -386 21 -384 24
rect -378 21 -376 24
rect -370 21 -368 24
rect -362 21 -360 24
rect -1189 -34 -1187 -31
rect -986 -40 -984 -37
rect -330 15 -328 18
rect -252 15 -250 18
rect -244 15 -242 18
rect -236 15 -234 18
rect -228 15 -226 18
rect -220 15 -218 18
rect -167 15 -165 18
rect -159 15 -157 18
rect -151 15 -149 18
rect -143 15 -141 18
rect -135 15 -133 18
rect -127 15 -125 18
rect -119 15 -117 18
rect -671 -26 -669 -23
rect -87 9 -85 12
rect -6 11 -4 14
rect 2 11 4 14
rect 10 11 12 14
rect 18 11 20 14
rect 26 11 28 14
rect 79 11 81 14
rect 87 11 89 14
rect 95 11 97 14
rect 103 11 105 14
rect 111 11 113 14
rect 119 11 121 14
rect 127 11 129 14
rect -418 -35 -416 -32
rect 159 5 161 8
rect -175 -41 -173 -38
rect 71 -45 73 -42
<< polycontact >>
rect -1558 12 -1554 16
rect -1614 -15 -1610 -11
rect -1304 16 -1300 20
rect -1646 -38 -1642 -34
rect -1360 -11 -1356 -7
rect -1105 9 -1101 13
rect -1392 -34 -1388 -30
rect -1466 -38 -1462 -34
rect -1434 -38 -1430 -34
rect -1161 -18 -1157 -14
rect -902 3 -898 7
rect -587 17 -583 21
rect -1267 -34 -1263 -30
rect -1235 -34 -1231 -30
rect -1193 -41 -1189 -37
rect -958 -24 -954 -20
rect -1064 -41 -1060 -37
rect -1032 -41 -1028 -37
rect -990 -47 -986 -43
rect -643 -10 -639 -6
rect -334 8 -330 12
rect -675 -33 -671 -29
rect -390 -19 -386 -15
rect -91 2 -87 6
rect -496 -33 -492 -29
rect -464 -33 -460 -29
rect -749 -47 -745 -43
rect -717 -47 -713 -43
rect -422 -42 -418 -38
rect -147 -25 -143 -21
rect 155 -2 159 2
rect -253 -42 -249 -38
rect -221 -42 -217 -38
rect -179 -48 -175 -44
rect 99 -29 103 -25
rect -7 -48 -3 -44
rect 25 -48 29 -44
rect 67 -52 71 -48
<< ndcontact >>
rect -1559 5 -1555 9
rect -1724 0 -1720 4
rect -1708 0 -1704 4
rect -1700 0 -1696 4
rect -1692 0 -1688 4
rect -1684 0 -1680 4
rect -1639 0 -1635 4
rect -1631 0 -1627 4
rect -1623 0 -1619 4
rect -1615 0 -1611 4
rect -1607 0 -1603 4
rect -1583 0 -1579 4
rect -1551 5 -1547 9
rect -1305 9 -1301 13
rect -1470 4 -1466 8
rect -1454 4 -1450 8
rect -1446 4 -1442 8
rect -1438 4 -1434 8
rect -1430 4 -1426 8
rect -1385 4 -1381 8
rect -1377 4 -1373 8
rect -1369 4 -1365 8
rect -1361 4 -1357 8
rect -1353 4 -1349 8
rect -1329 4 -1325 8
rect -1297 9 -1293 13
rect -1106 2 -1102 6
rect -1271 -3 -1267 1
rect -1255 -3 -1251 1
rect -1247 -3 -1243 1
rect -1239 -3 -1235 1
rect -1231 -3 -1227 1
rect -1186 -3 -1182 1
rect -1178 -3 -1174 1
rect -1170 -3 -1166 1
rect -1162 -3 -1158 1
rect -1154 -3 -1150 1
rect -1130 -3 -1126 1
rect -1098 2 -1094 6
rect -588 10 -584 14
rect -753 5 -749 9
rect -903 -4 -899 0
rect -1068 -9 -1064 -5
rect -1393 -41 -1389 -37
rect -1647 -45 -1643 -41
rect -1639 -45 -1635 -41
rect -1385 -41 -1381 -37
rect -1052 -9 -1048 -5
rect -1044 -9 -1040 -5
rect -1036 -9 -1032 -5
rect -1028 -9 -1024 -5
rect -983 -9 -979 -5
rect -975 -9 -971 -5
rect -967 -9 -963 -5
rect -959 -9 -955 -5
rect -951 -9 -947 -5
rect -927 -9 -923 -5
rect -895 -4 -891 0
rect -1194 -48 -1190 -44
rect -1186 -48 -1182 -44
rect -737 5 -733 9
rect -729 5 -725 9
rect -721 5 -717 9
rect -713 5 -709 9
rect -668 5 -664 9
rect -660 5 -656 9
rect -652 5 -648 9
rect -644 5 -640 9
rect -636 5 -632 9
rect -612 5 -608 9
rect -580 10 -576 14
rect -335 1 -331 5
rect -500 -4 -496 0
rect -484 -4 -480 0
rect -476 -4 -472 0
rect -468 -4 -464 0
rect -460 -4 -456 0
rect -415 -4 -411 0
rect -407 -4 -403 0
rect -399 -4 -395 0
rect -391 -4 -387 0
rect -383 -4 -379 0
rect -359 -4 -355 0
rect -327 1 -323 5
rect -92 -5 -88 -1
rect -257 -10 -253 -6
rect -676 -40 -672 -36
rect -668 -40 -664 -36
rect -241 -10 -237 -6
rect -233 -10 -229 -6
rect -225 -10 -221 -6
rect -217 -10 -213 -6
rect -172 -10 -168 -6
rect -164 -10 -160 -6
rect -156 -10 -152 -6
rect -148 -10 -144 -6
rect -140 -10 -136 -6
rect -116 -10 -112 -6
rect -84 -5 -80 -1
rect 154 -9 158 -5
rect -11 -14 -7 -10
rect -423 -49 -419 -45
rect -991 -54 -987 -50
rect -983 -54 -979 -50
rect -415 -49 -411 -45
rect 5 -14 9 -10
rect 13 -14 17 -10
rect 21 -14 25 -10
rect 29 -14 33 -10
rect 74 -14 78 -10
rect 82 -14 86 -10
rect 90 -14 94 -10
rect 98 -14 102 -10
rect 106 -14 110 -10
rect 130 -14 134 -10
rect 162 -9 166 -5
rect -180 -55 -176 -51
rect -172 -55 -168 -51
rect 66 -59 70 -55
rect 74 -59 78 -55
<< pdcontact >>
rect -1724 25 -1720 29
rect -1716 25 -1712 29
rect -1708 25 -1704 29
rect -1700 25 -1696 29
rect -1684 25 -1680 29
rect -1639 25 -1635 29
rect -1615 25 -1611 29
rect -1607 25 -1603 29
rect -1599 25 -1595 29
rect -1591 25 -1587 29
rect -1583 25 -1579 29
rect -1470 29 -1466 33
rect -1462 29 -1458 33
rect -1454 29 -1450 33
rect -1446 29 -1442 33
rect -1430 29 -1426 33
rect -1385 29 -1381 33
rect -1361 29 -1357 33
rect -1353 29 -1349 33
rect -1345 29 -1341 33
rect -1337 29 -1333 33
rect -1329 29 -1325 33
rect -1559 19 -1555 23
rect -1551 19 -1547 23
rect -1305 23 -1301 27
rect -1297 23 -1293 27
rect -1271 22 -1267 26
rect -1263 22 -1259 26
rect -1255 22 -1251 26
rect -1247 22 -1243 26
rect -1231 22 -1227 26
rect -1186 22 -1182 26
rect -1162 22 -1158 26
rect -1154 22 -1150 26
rect -1146 22 -1142 26
rect -1138 22 -1134 26
rect -753 30 -749 34
rect -745 30 -741 34
rect -737 30 -733 34
rect -729 30 -725 34
rect -713 30 -709 34
rect -668 30 -664 34
rect -644 30 -640 34
rect -636 30 -632 34
rect -628 30 -624 34
rect -620 30 -616 34
rect -612 30 -608 34
rect -1130 22 -1126 26
rect -1647 -31 -1643 -27
rect -1639 -31 -1635 -27
rect -1106 16 -1102 20
rect -1098 16 -1094 20
rect -1068 16 -1064 20
rect -1060 16 -1056 20
rect -1052 16 -1048 20
rect -1044 16 -1040 20
rect -1028 16 -1024 20
rect -983 16 -979 20
rect -959 16 -955 20
rect -951 16 -947 20
rect -943 16 -939 20
rect -935 16 -931 20
rect -927 16 -923 20
rect -1393 -27 -1389 -23
rect -1385 -27 -1381 -23
rect -903 10 -899 14
rect -895 10 -891 14
rect -588 24 -584 28
rect -580 24 -576 28
rect -500 21 -496 25
rect -492 21 -488 25
rect -484 21 -480 25
rect -476 21 -472 25
rect -460 21 -456 25
rect -415 21 -411 25
rect -391 21 -387 25
rect -383 21 -379 25
rect -375 21 -371 25
rect -367 21 -363 25
rect -359 21 -355 25
rect -1194 -34 -1190 -30
rect -1186 -34 -1182 -30
rect -991 -40 -987 -36
rect -983 -40 -979 -36
rect -335 15 -331 19
rect -327 15 -323 19
rect -257 15 -253 19
rect -249 15 -245 19
rect -241 15 -237 19
rect -233 15 -229 19
rect -217 15 -213 19
rect -172 15 -168 19
rect -148 15 -144 19
rect -140 15 -136 19
rect -132 15 -128 19
rect -124 15 -120 19
rect -116 15 -112 19
rect -676 -26 -672 -22
rect -668 -26 -664 -22
rect -92 9 -88 13
rect -84 9 -80 13
rect -11 11 -7 15
rect -3 11 1 15
rect 5 11 9 15
rect 13 11 17 15
rect 29 11 33 15
rect 74 11 78 15
rect 98 11 102 15
rect 106 11 110 15
rect 114 11 118 15
rect 122 11 126 15
rect 130 11 134 15
rect -423 -35 -419 -31
rect -415 -35 -411 -31
rect 154 5 158 9
rect 162 5 166 9
rect -180 -41 -176 -37
rect -172 -41 -168 -37
rect 66 -45 70 -41
rect 74 -45 78 -41
<< psubstratepcontact >>
rect -1725 -8 -1721 -4
rect -1692 -8 -1688 -4
rect -1640 -8 -1636 -4
rect -1623 -8 -1619 -4
rect -1559 -3 -1555 1
rect -1471 -4 -1467 0
rect -1582 -8 -1578 -4
rect -1438 -4 -1434 0
rect -1386 -4 -1382 0
rect -1369 -4 -1365 0
rect -1305 1 -1301 5
rect -1328 -4 -1324 0
rect -1272 -11 -1268 -7
rect -1239 -11 -1235 -7
rect -1187 -11 -1183 -7
rect -1170 -11 -1166 -7
rect -1106 -6 -1102 -2
rect -1129 -11 -1125 -7
rect -1069 -17 -1065 -13
rect -1647 -53 -1643 -49
rect -1393 -49 -1389 -45
rect -1036 -17 -1032 -13
rect -984 -17 -980 -13
rect -967 -17 -963 -13
rect -903 -12 -899 -8
rect -754 -3 -750 1
rect -926 -17 -922 -13
rect -1194 -56 -1190 -52
rect -721 -3 -717 1
rect -669 -3 -665 1
rect -652 -3 -648 1
rect -588 2 -584 6
rect -611 -3 -607 1
rect -501 -12 -497 -8
rect -468 -12 -464 -8
rect -416 -12 -412 -8
rect -399 -12 -395 -8
rect -335 -7 -331 -3
rect -358 -12 -354 -8
rect -258 -18 -254 -14
rect -676 -48 -672 -44
rect -225 -18 -221 -14
rect -173 -18 -169 -14
rect -156 -18 -152 -14
rect -92 -13 -88 -9
rect -115 -18 -111 -14
rect -12 -22 -8 -18
rect -991 -62 -987 -58
rect -423 -57 -419 -53
rect 21 -22 25 -18
rect 73 -22 77 -18
rect 90 -22 94 -18
rect 154 -17 158 -13
rect 131 -22 135 -18
rect -180 -63 -176 -59
rect 66 -67 70 -63
<< nsubstratencontact >>
rect -1446 42 -1442 46
rect -1700 38 -1696 42
rect -1361 41 -1357 45
rect -729 43 -725 47
rect -644 42 -640 46
rect -1615 37 -1611 41
rect -1559 27 -1555 31
rect -1247 35 -1243 39
rect -1305 31 -1301 35
rect -1162 34 -1158 38
rect -1044 29 -1040 33
rect -959 28 -955 32
rect -588 32 -584 36
rect -476 34 -472 38
rect -391 33 -387 37
rect -1106 24 -1102 28
rect -1647 -23 -1643 -19
rect -903 18 -899 22
rect -1393 -19 -1389 -15
rect -233 28 -229 32
rect -148 27 -144 31
rect -335 23 -331 27
rect -1194 -26 -1190 -22
rect -991 -32 -987 -28
rect 13 24 17 28
rect 98 23 102 27
rect -92 17 -88 21
rect -676 -18 -672 -14
rect 154 13 158 17
rect -423 -27 -419 -23
rect -180 -33 -176 -29
rect 66 -37 70 -33
<< labels >>
rlabel metal1 -13 24 35 27 1 VDD
rlabel metal1 -13 -22 35 -19 5 GND
rlabel polysilicon 18 -10 20 11 0 B
rlabel polysilicon 26 -10 28 11 0 Cin
rlabel metal1 -13 -1 35 2 3 Cout'
rlabel metal1 72 24 136 27 1 VDD
rlabel metal1 72 -22 136 -19 5 GND
rlabel polysilicon 119 -10 121 11 0 B
rlabel polysilicon 127 -10 129 11 0 Cin
rlabel metal1 75 -51 86 -48 3 Cout
rlabel metal1 66 -37 78 -34 1 VDD
rlabel metal1 66 -66 78 -63 5 GND
rlabel metal1 154 13 166 16 1 VDD
rlabel metal1 154 -16 166 -13 5 GND
rlabel metal1 72 -1 155 2 1 Sout'
rlabel metal1 163 -1 175 2 3 Sout
rlabel polysilicon 111 -10 113 11 0 A
rlabel polysilicon 95 -10 97 11 0 Cin
rlabel polysilicon 87 -10 89 11 0 B
rlabel polysilicon 79 -10 81 11 0 A
rlabel polysilicon 10 -10 12 11 0 A
rlabel polysilicon -6 -10 -4 11 0 Cin
rlabel metal1 -83 3 -71 6 3 Sout
rlabel metal1 -174 3 -91 6 1 Sout'
rlabel metal1 -92 -12 -80 -9 5 GND
rlabel metal1 -92 17 -80 20 1 VDD
rlabel metal1 -180 -62 -168 -59 5 GND
rlabel metal1 -180 -33 -168 -30 1 VDD
rlabel metal1 -171 -47 -160 -44 3 Cout
rlabel polysilicon -167 -6 -165 15 0 A
rlabel metal1 -174 -18 -110 -15 5 GND
rlabel metal1 -174 28 -110 31 1 VDD
rlabel metal1 -259 3 -211 6 3 Cout'
rlabel polysilicon -220 -6 -218 15 0 Cin
rlabel polysilicon -228 -6 -226 15 0 B
rlabel polysilicon -236 -6 -234 15 0 A
rlabel polysilicon -244 -6 -242 15 0 B
rlabel polysilicon -252 -6 -250 15 0 Cin
rlabel metal1 -259 -18 -211 -15 5 GND
rlabel metal1 -259 28 -211 31 1 VDD
rlabel metal1 -326 9 -314 12 3 Sout
rlabel metal1 -417 9 -334 12 1 Sout'
rlabel metal1 -335 -6 -323 -3 5 GND
rlabel metal1 -335 23 -323 26 1 VDD
rlabel metal1 -423 -56 -411 -53 5 GND
rlabel metal1 -423 -27 -411 -24 1 VDD
rlabel metal1 -414 -41 -403 -38 3 Cout
rlabel polysilicon -362 0 -360 21 0 Cin
rlabel polysilicon -370 0 -368 21 0 B
rlabel polysilicon -378 0 -376 21 0 A
rlabel polysilicon -394 0 -392 21 0 Cin
rlabel polysilicon -402 0 -400 21 0 B
rlabel polysilicon -410 0 -408 21 0 A
rlabel metal1 -417 -12 -353 -9 5 GND
rlabel metal1 -417 34 -353 37 1 VDD
rlabel metal1 -502 9 -454 12 3 Cout'
rlabel polysilicon -463 0 -461 21 0 Cin
rlabel polysilicon -471 0 -469 21 0 B
rlabel polysilicon -479 0 -477 21 0 A
rlabel polysilicon -487 0 -485 21 0 B
rlabel polysilicon -495 0 -493 21 0 Cin
rlabel metal1 -502 -12 -454 -9 5 GND
rlabel metal1 -502 34 -454 37 1 VDD
rlabel polysilicon -159 -6 -157 15 0 B
rlabel polysilicon -151 -6 -149 15 0 Cin
rlabel polysilicon -135 -6 -133 15 0 A
rlabel polysilicon -127 -6 -125 15 0 B
rlabel polysilicon -119 -6 -117 15 0 Cin
rlabel polysilicon 2 -10 4 11 0 B
rlabel metal1 -755 43 -707 46 1 VDD
rlabel metal1 -755 -3 -707 0 5 GND
rlabel polysilicon -748 9 -746 30 0 Cin
rlabel polysilicon -740 9 -738 30 0 B
rlabel polysilicon -732 9 -730 30 0 A
rlabel polysilicon -724 9 -722 30 0 B
rlabel polysilicon -716 9 -714 30 0 Cin
rlabel metal1 -755 18 -707 21 3 Cout'
rlabel metal1 -670 43 -606 46 1 VDD
rlabel metal1 -670 -3 -606 0 5 GND
rlabel polysilicon -663 9 -661 30 0 A
rlabel polysilicon -655 9 -653 30 0 B
rlabel polysilicon -647 9 -645 30 0 Cin
rlabel polysilicon -631 9 -629 30 0 A
rlabel polysilicon -623 9 -621 30 0 B
rlabel polysilicon -615 9 -613 30 0 Cin
rlabel metal1 -667 -32 -656 -29 3 Cout
rlabel metal1 -676 -18 -664 -15 1 VDD
rlabel metal1 -676 -47 -664 -44 5 GND
rlabel metal1 -588 32 -576 35 1 VDD
rlabel metal1 -588 3 -576 6 5 GND
rlabel metal1 -670 18 -587 21 1 Sout'
rlabel metal1 -579 18 -567 21 3 Sout
rlabel metal1 -1070 29 -1022 32 1 VDD
rlabel metal1 -1070 -17 -1022 -14 5 GND
rlabel polysilicon -1063 -5 -1061 16 0 Cin
rlabel polysilicon -1055 -5 -1053 16 0 B
rlabel polysilicon -1047 -5 -1045 16 0 A
rlabel polysilicon -1039 -5 -1037 16 0 B
rlabel polysilicon -1031 -5 -1029 16 0 Cin
rlabel metal1 -1070 4 -1022 7 3 Cout'
rlabel metal1 -985 29 -921 32 1 VDD
rlabel metal1 -985 -17 -921 -14 5 GND
rlabel polysilicon -978 -5 -976 16 0 A
rlabel polysilicon -970 -5 -968 16 0 B
rlabel polysilicon -962 -5 -960 16 0 Cin
rlabel polysilicon -946 -5 -944 16 0 A
rlabel polysilicon -938 -5 -936 16 0 B
rlabel polysilicon -930 -5 -928 16 0 Cin
rlabel metal1 -982 -46 -971 -43 3 Cout
rlabel metal1 -991 -32 -979 -29 1 VDD
rlabel metal1 -991 -61 -979 -58 5 GND
rlabel metal1 -903 18 -891 21 1 VDD
rlabel metal1 -903 -11 -891 -8 5 GND
rlabel metal1 -985 4 -902 7 1 Sout'
rlabel metal1 -894 4 -882 7 3 Sout
rlabel metal1 -1296 17 -1284 20 3 Sout
rlabel metal1 -1387 17 -1304 20 1 Sout'
rlabel metal1 -1305 2 -1293 5 5 GND
rlabel metal1 -1305 31 -1293 34 1 VDD
rlabel metal1 -1393 -48 -1381 -45 5 GND
rlabel metal1 -1393 -19 -1381 -16 1 VDD
rlabel metal1 -1384 -33 -1373 -30 3 Cout
rlabel polysilicon -1332 8 -1330 29 0 Cin
rlabel polysilicon -1340 8 -1338 29 0 B
rlabel polysilicon -1348 8 -1346 29 0 A
rlabel polysilicon -1364 8 -1362 29 0 Cin
rlabel polysilicon -1372 8 -1370 29 0 B
rlabel polysilicon -1380 8 -1378 29 0 A
rlabel metal1 -1387 -4 -1323 -1 5 GND
rlabel metal1 -1387 42 -1323 45 1 VDD
rlabel metal1 -1472 17 -1424 20 3 Cout'
rlabel polysilicon -1433 8 -1431 29 0 Cin
rlabel polysilicon -1441 8 -1439 29 0 B
rlabel polysilicon -1449 8 -1447 29 0 A
rlabel polysilicon -1457 8 -1455 29 0 B
rlabel polysilicon -1465 8 -1463 29 0 Cin
rlabel metal1 -1472 -4 -1424 -1 5 GND
rlabel metal1 -1472 42 -1424 45 1 VDD
rlabel polysilicon -1258 1 -1256 22 0 B
rlabel polysilicon -1266 1 -1264 22 0 Cin
rlabel polysilicon -1250 1 -1248 22 0 A
rlabel polysilicon -1181 1 -1179 22 0 A
rlabel polysilicon -1173 1 -1171 22 0 B
rlabel polysilicon -1165 1 -1163 22 0 Cin
rlabel polysilicon -1149 1 -1147 22 0 A
rlabel metal1 -1097 10 -1085 13 3 Sout
rlabel metal1 -1188 10 -1105 13 1 Sout'
rlabel metal1 -1106 -5 -1094 -2 5 GND
rlabel metal1 -1106 24 -1094 27 1 VDD
rlabel metal1 -1194 -55 -1182 -52 5 GND
rlabel metal1 -1194 -26 -1182 -23 1 VDD
rlabel metal1 -1185 -40 -1174 -37 3 Cout
rlabel polysilicon -1133 1 -1131 22 0 Cin
rlabel polysilicon -1141 1 -1139 22 0 B
rlabel metal1 -1188 -11 -1124 -8 5 GND
rlabel metal1 -1188 35 -1124 38 1 VDD
rlabel metal1 -1273 10 -1225 13 3 Cout'
rlabel polysilicon -1234 1 -1232 22 0 Cin
rlabel polysilicon -1242 1 -1240 22 0 B
rlabel metal1 -1273 -11 -1225 -8 5 GND
rlabel metal1 -1273 35 -1225 38 1 VDD
rlabel polysilicon -1711 4 -1709 25 0 B
rlabel polysilicon -1719 4 -1717 25 0 Cin
rlabel polysilicon -1703 4 -1701 25 0 A
rlabel polysilicon -1634 4 -1632 25 0 A
rlabel polysilicon -1626 4 -1624 25 0 B
rlabel polysilicon -1618 4 -1616 25 0 Cin
rlabel polysilicon -1602 4 -1600 25 0 A
rlabel metal1 -1550 13 -1538 16 3 Sout
rlabel metal1 -1641 13 -1558 16 1 Sout'
rlabel metal1 -1559 -2 -1547 1 5 GND
rlabel metal1 -1559 27 -1547 30 1 VDD
rlabel metal1 -1647 -52 -1635 -49 5 GND
rlabel metal1 -1647 -23 -1635 -20 1 VDD
rlabel metal1 -1638 -37 -1627 -34 3 Cout
rlabel polysilicon -1586 4 -1584 25 0 Cin
rlabel polysilicon -1594 4 -1592 25 0 B
rlabel metal1 -1641 -8 -1577 -5 5 GND
rlabel metal1 -1641 38 -1577 41 1 VDD
rlabel metal1 -1726 13 -1678 16 3 Cout'
rlabel polysilicon -1687 4 -1685 25 0 Cin
rlabel polysilicon -1695 4 -1693 25 0 B
rlabel metal1 -1726 -8 -1678 -5 5 GND
rlabel metal1 -1726 38 -1678 41 1 VDD
<< end >>
